module c5315(G1,G4,G11,G14,G17,G20,G23,G24,G25,G26,G27,
      G31,G34,G37,G40,G43,G46,G49,G52,G53,G54,G61,
      G64,G67,G70,G73,G76,G79,G80,G81,G82,G83,G86,
      G87,G88,G91,G94,G97,G100,G103,G106,G109,G112,G113,
      G114,G115,G116,G117,G118,G119,G120,G121,G122,G123,G126,
      G127,G128,G129,G130,G131,G132,G135,G136,G137,G140,G141,
      G145,G146,G149,G152,G155,G158,G161,G164,G167,G170,G173,
      G176,G179,G182,G185,G188,G191,G194,G197,G200,G203,G206,
      G209,G210,G217,G218,G225,G226,G233,G234,G241,G242,G245,
      G248,G251,G254,G257,G264,G265,G272,G273,G280,G281,G288,
      G289,G292,G293,G299,G302,G307,G308,G315,G316,G323,G324,
      G331,G332,G335,G338,G341,G348,G351,G358,G361,G366,G369,
      G372,G373,G374,G386,G389,G400,G411,G422,G435,G446,G457,
      G468,G479,G490,G503,G514,G523,G534,G545,G549,G552,G556,
      G559,G562,G1497,G1689,G1690,G1691,G1694,G2174,G2358,G2824,G3173,
      G3546,G3548,G3550,G3552,G3717,G3724,G4087,G4088,G4089,G4090,G4091,
      G4092,G4115,G144,G298,G973,G594,G599,G600,G601,G602,G603,
      G604,G611,G612,G810,G848,G849,G850,G851,G634,G815,G845,
      G847,G926,G923,G921,G892,G887,G606,G656,G809,G993,G978,
      G949,G939,G889,G593,G636,G704,G717,G820,G639,G673,G707,
      G715,G598,G610,G588,G615,G626,G632,G1002,G1004,G591,G618,
      G621,G629,G822,G838,G861,G623,G722,G832,G834,G836,G859,
      G871,G873,G875,G877,G998,G1000,G575,G585,G661,G693,G747,
      G752,G757,G762,G787,G792,G797,G802,G642,G664,G667,G670,
      G676,G696,G699,G702,G818,G813,G824,G826,G828,G830,G854,
      G863,G865,G867,G869,G712,G727,G732,G737,G742,G772,G777,
      G782,G645,G648,G651,G654,G679,G682,G685,G688,G843,G882,
      G767,G807,G658,G690);

input G1,G4,G11,G14,G17,G20,G23,G24,G25,G26,G27,
      G31,G34,G37,G40,G43,G46,G49,G52,G53,G54,G61,
      G64,G67,G70,G73,G76,G79,G80,G81,G82,G83,G86,
      G87,G88,G91,G94,G97,G100,G103,G106,G109,G112,G113,
      G114,G115,G116,G117,G118,G119,G120,G121,G122,G123,G126,
      G127,G128,G129,G130,G131,G132,G135,G136,G137,G140,G141,
      G145,G146,G149,G152,G155,G158,G161,G164,G167,G170,G173,
      G176,G179,G182,G185,G188,G191,G194,G197,G200,G203,G206,
      G209,G210,G217,G218,G225,G226,G233,G234,G241,G242,G245,
      G248,G251,G254,G257,G264,G265,G272,G273,G280,G281,G288,
      G289,G292,G293,G299,G302,G307,G308,G315,G316,G323,G324,
      G331,G332,G335,G338,G341,G348,G351,G358,G361,G366,G369,
      G372,G373,G374,G386,G389,G400,G411,G422,G435,G446,G457,
      G468,G479,G490,G503,G514,G523,G534,G545,G549,G552,G556,
      G559,G562,G1497,G1689,G1690,G1691,G1694,G2174,G2358,G2824,G3173,
      G3546,G3548,G3550,G3552,G3717,G3724,G4087,G4088,G4089,G4090,G4091,
      G4092,G4115;

output G144,G298,G973,G594,G599,G600,G601,G602,G603,G604,G611,
       G612,G810,G848,G849,G850,G851,G634,G815,G845,G847,G926,
       G923,G921,G892,G887,G606,G656,G809,G993,G978,G949,G939,
       G889,G593,G636,G704,G717,G820,G639,G673,G707,G715,G598,
       G610,G588,G615,G626,G632,G1002,G1004,G591,G618,G621,G629,
       G822,G838,G861,G623,G722,G832,G834,G836,G859,G871,G873,
       G875,G877,G998,G1000,G575,G585,G661,G693,G747,G752,G757,
       G762,G787,G792,G797,G802,G642,G664,G667,G670,G676,G696,
       G699,G702,G818,G813,G824,G826,G828,G830,G854,G863,G865,
       G867,G869,G712,G727,G732,G737,G742,G772,G777,G782,G645,
       G648,G651,G654,G679,G682,G685,G688,G843,G882,G767,G807,
       G658,G690;

wire G4114,G2825,G3547,G3549,G3551,G3553,G633,G814,G816,G844,G846,
     G852,G1502,G1528,G1552,G1609,G1633,G1697,G1698,G1701,G2179,G2203,
     G2226,G2281,G2304,G2361,G2370,G2382,G2393,G2405,G2418,G2442,G2476,
     G2500,G2533,G2537,G2541,G2545,G2549,G2553,G2557,G2561,G2627,G2631,
     G2635,G2639,G2643,G2647,G2651,G2655,G2721,G2734,G2816,G2822,G2826,
     G2828,G2882,G2886,G2890,G2894,G2898,G2902,G2948,G2952,G2956,G2960,
     G2964,G2968,G3024,G3028,G3032,G3036,G3040,G3044,G3048,G3052,G3092,
     G3105,G3175,G3176,G3181,G3204,G3208,G3212,G3216,G3220,G3224,G3256,
     G3260,G3264,G3268,G3272,G3276,G3302,G3314,G3354,G3358,G3362,G3366,
     G3370,G3374,G3378,G3382,G3440,G3554,G3555,G3556,G3558,G3582,G3616,
     G3628,G3660,G3684,G3721,G3728,G3737,G3757,G3795,G3815,G3972,G3991,
     G4030,G4049,G4110,G4119,G4127,G4135,G4143,G4151,G4159,G4167,G4175,
     G4183,G4188,G4276,G4284,G4292,G4300,G4308,G4316,G4324,G4332,G4340,
     G4631,G4639,G4647,G4655,G4663,G4671,G4676,G4764,G4772,G4780,G4788,
     G4796,G4804,G5082,G5085,G5090,G5093,G5098,G5101,G5108,G5111,G5332,
     G5335,G5340,G5343,G5348,G5351,G5356,G5359,G5369,G2979,G2999,G1580,
     G1586,G1592,G1598,G1604,G1668,G1674,G1680,G1686,G2254,G2260,G2266,
     G2272,G2278,G2339,G2345,G2351,G2357,G711,G721,G726,G731,G736,
     G741,G746,G751,G756,G761,G766,G771,G776,G781,G786,G791,
     G796,G801,G806,G3734,G842,G858,G881,G4123,G4131,G4139,G4147,
     G4155,G4163,G4171,G4179,G4187,G4194,G4282,G4290,G4298,G4306,G4314,
     G4322,G4330,G4338,G4346,G1526,G1540,G1564,G1606,G1621,G1645,G1661,
     G1688,G4635,G4643,G4651,G4659,G4667,G4675,G4682,G4770,G4778,G4786,
     G4794,G4802,G4810,G2202,G2215,G2238,G2279,G2293,G2316,G2332,G2430,
     G2454,G2488,G2512,G2536,G2540,G2544,G2548,G2552,G2556,G2560,G2564,
     G2566,G2572,G2578,G2584,G2590,G2595,G2600,G2605,G2630,G2634,G2638,
     G2642,G2646,G2650,G2654,G2658,G2660,G2666,G2672,G2678,G2684,G2689,
     G2694,G2699,G2728,G2741,G2748,G2750,G2752,G2754,G2756,G2758,G2760,
     G2762,G2764,G2766,G2827,G2838,G2847,G2885,G2889,G2893,G2897,G2901,
     G2905,G2906,G2909,G2913,G2918,G2922,G2927,G2951,G2955,G2959,G2963,
     G2967,G2971,G2973,G2980,G2982,G2988,G2994,G3001,G3006,G3027,G3031,
     G3035,G3039,G3043,G3047,G3051,G3055,G3056,G3060,G3064,G3068,G3073,
     G3078,G3083,G3088,G3099,G3112,G3119,G3121,G3123,G3125,G3126,G3128,
     G3130,G3132,G3134,G3136,G3187,G3193,G3196,G3199,G3202,G3207,G3211,
     G3215,G3219,G3223,G3227,G3228,G3232,G3234,G3238,G3243,G3247,G3249,
     G3253,G3259,G3263,G3267,G3271,G3275,G3279,G3280,G3283,G3287,G3292,
     G3295,G3299,G3305,G3306,G3310,G3317,G3318,G3322,G3326,G3333,G3357,
     G3361,G3365,G3369,G3373,G3377,G3381,G3385,G3386,G3390,G3394,G3398,
     G3403,G3408,G3413,G3418,G5088,G5089,G5096,G5097,G3489,G3493,G3570,
     G3594,G3622,G3632,G3637,G3640,G3643,G3646,G3672,G3696,G3745,G3765,
     G3803,G3823,G5338,G5339,G5346,G5347,G5354,G5355,G3979,G3998,G4037,
     G4056,G4094,G5104,G5105,G5114,G5115,G5362,G5363,G5366,G5373,G2568,
     G2574,G2580,G2586,G2592,G2597,G2602,G2607,G2662,G2668,G2674,G2680,
     G2686,G2691,G2696,G2701,G2907,G2910,G2914,G2920,G2924,G2929,G2975,
     G2984,G2990,G2996,G3003,G3008,G3015,G3057,G3061,G3065,G3069,G3075,
     G3080,G3085,G3090,G3229,G3233,G3235,G3239,G3244,G3250,G3254,G3281,
     G3284,G3288,G3293,G3296,G3300,G3327,G3334,G3387,G3391,G3395,G3399,
     G3405,G3410,G3415,G3420,G3422,G3423,G3431,G3432,G3895,G3896,G3904,
     G3905,G3913,G3914,G5106,G5107,G5116,G5117,G5364,G5365,G2880,G2881,
     G1579,G1585,G1591,G1597,G1603,G1667,G1673,G1679,G1685,G2876,G2877,
     G2253,G2259,G2265,G2271,G2277,G2338,G2344,G2350,G2356,G2868,G2869,
     G710,G2872,G2873,G720,G725,G730,G735,G740,G745,G750,G755,
     G760,G765,G770,G775,G780,G785,G790,G795,G800,G805,G841,
     G857,G880,G1660,G2331,G2569,G2575,G2581,G2587,G2593,G2598,G2603,
     G2608,G2663,G2669,G2675,G2681,G2687,G2692,G2697,G2702,G2747,G2749,
     G2751,G2753,G2755,G2757,G2759,G2761,G2763,G2765,G2857,G2908,G2911,
     G2915,G2925,G2930,G2933,G2976,G2985,G2991,G2997,G3004,G3009,G3058,
     G3062,G3066,G3070,G3076,G3081,G3086,G3091,G3118,G3120,G3122,G3124,
     G3127,G3129,G3131,G3133,G3135,G3147,G3192,G3195,G3198,G3201,G3230,
     G3236,G3240,G3245,G3251,G3255,G3282,G3285,G3289,G3297,G3301,G3309,
     G3313,G3321,G3325,G3328,G3329,G3335,G3336,G3341,G3345,G3388,G3392,
     G3396,G3400,G3406,G3411,G3416,G3421,G3424,G3433,G3492,G3496,G3780,
     G3783,G3786,G3789,G3838,G3841,G3844,G3847,G3897,G3906,G3915,G4011,
     G4014,G4017,G4020,G4023,G4069,G4072,G4075,G4078,G4081,G5206,G5209,
     G5307,G5322,G5372,G5375,G5399,G2813,G3197,G3200,G3203,G3194,G2570,
     G2576,G2582,G2588,G2664,G2670,G2676,G2682,G2767,G2772,G2776,G2780,
     G2784,G2788,G2794,G2798,G2802,G2912,G2916,G2936,G2977,G2986,G2992,
     G3059,G3063,G3067,G3071,G3137,G3139,G3143,G3151,G3155,G3161,G3165,
     G3167,G3231,G3237,G3241,G3286,G3290,G3330,G3337,G3342,G3346,G3348,
     G3352,G3389,G3393,G3397,G3401,G3845,G5126,G5178,G5325,G5374,G2810,
     G635,G2878,G2879,G2874,G2875,G703,G2866,G2867,G2870,G2871,G716,
     G819,G1789,G2036,G2611,G2615,G2619,G2623,G2705,G2709,G2713,G2717,
     G2939,G2942,G2945,G3012,G3018,G3021,G3331,G3338,G3343,G3347,G3428,
     G3437,G3514,G3836,G3852,G5311,G3901,G3910,G3934,G3938,G4652,G4783,
     G5137,G5212,G5213,G5260,G5263,G5268,G5271,G5276,G5279,G5289,G5296,
     G5299,G5304,G5312,G5315,G5328,G5396,G5403,G1286,G2809,G597,G1031,
     G637,G671,G705,G713,G1046,G1064,G1071,G1097,G1111,G1128,G1145,
     G1160,G1301,G1318,G1324,G1341,G1359,G1382,G1404,G1412,G1704,G1712,
     G1724,G1742,G1749,G1775,G1806,G1823,G1829,G1837,G1958,G1966,G1978,
     G1995,G2001,G2018,G2059,G2081,G2089,G2106,G3170,G3332,G3339,G5132,
     G5184,G3853,G3874,G4076,G4116,G4124,G4132,G4140,G4148,G4156,G4164,
     G4172,G4180,G4228,G4279,G4287,G4295,G4303,G4311,G4319,G4327,G4335,
     G4343,G4348,G4464,G4628,G4636,G4644,G4660,G4668,G4716,G4767,G4775,
     G4791,G4799,G4807,G4812,G5118,G5121,G5129,G5134,G5142,G5145,G5152,
     G5155,G5162,G5165,G5170,G5173,G5181,G5186,G5189,G5196,G5199,G5214,
     G5215,G5329,G5330,G2807,G2808,G2811,G2812,G2814,G2626,G2622,G2618,
     G2614,G2720,G2716,G2712,G2708,G3731,G4658,G1777,G2019,G4787,G3350,
     G3353,G5141,G3513,G3516,G3517,G3778,G3781,G3784,G3787,G3839,G3842,
     G5266,G5267,G5274,G5275,G5302,G5303,G5310,G3891,G3937,G3941,G3955,
     G3958,G4009,G4012,G4015,G4018,G4067,G4070,G4073,G4079,G5239,G5282,
     G5283,G5293,G5318,G5319,G5331,G5402,G5405,G595,G596,G607,G608,
     G1845,G1846,G2115,G2116,G4122,G1022,G4130,G1033,G4138,G1051,G4146,
     G1079,G4154,G1088,G4162,G1099,G4170,G1115,G4178,G1133,G4186,G1151,
     G4234,G1276,G4283,G1287,G4291,G1305,G4299,G1330,G4307,G1342,G4315,
     G1363,G4323,G1388,G4331,G1420,G4339,G1428,G4347,G4634,G1729,G4642,
     G1757,G4650,G1766,G1776,G4666,G1793,G4674,G1811,G1849,G1852,G1875,
     G4722,G1982,G4771,G2007,G4779,G2020,G2040,G4795,G2065,G4803,G2097,
     G4811,G2119,G2122,G5124,G5125,G3452,G5133,G5140,G3462,G5168,G5169,
     G5176,G5177,G3484,G5185,G3515,G3518,G3857,G3860,G3861,G3869,G3870,
     G3878,G3881,G3882,G3890,G3954,G3957,G4021,G4099,G4236,G4354,G4406,
     G4470,G4552,G4679,G4687,G4695,G4703,G4711,G4724,G4818,G4855,G4865,
     G4870,G4913,G4923,G4951,G5006,G5039,G5148,G5149,G5158,G5159,G5192,
     G5193,G5202,G5203,G5284,G5285,G5320,G5321,G5386,G5404,G609,G1021,
     G1032,G1050,G1078,G1087,G1098,G1114,G1132,G1150,G1277,G1288,G1306,
     G1331,G1343,G1364,G1389,G1421,G1429,G1728,G1756,G1765,G1778,G1792,
     G1810,G1983,G2008,G2021,G2041,G2066,G2098,G3443,G3444,G3453,G3461,
     G3466,G3467,G3475,G3476,G3485,G5243,G3862,G3871,G3883,G3892,G3956,
     G3959,G4756,G5150,G5151,G5160,G5161,G5194,G5195,G5204,G5205,G5236,
     G5286,G5379,G5389,G5425,G1023,G1034,G1052,G1080,G1089,G1100,G1116,
     G1134,G1152,G4242,G1278,G1289,G1307,G1332,G1344,G1365,G1390,G1422,
     G1430,G1730,G1758,G1767,G1794,G1812,G1876,G4683,G4691,G4699,G4707,
     G4715,G4730,G1984,G2009,G2042,G2067,G2099,G4869,G4927,G3445,G3454,
     G3463,G3468,G3477,G3486,G4103,G4412,G4558,G4859,G4876,G4917,G4955,
     G5012,G5043,G5216,G5219,G5226,G5229,G5392,G5422,G1866,G1877,G4762,
     G2142,G2146,G5242,G3532,G3866,G3887,G3918,G3922,G3926,G3930,G5429,
     G4104,G4743,G4991,G5001,G5292,G5295,G5383,G5393,G5394,G1439,G1440,
     G1441,G1847,G1168,G1169,G1170,G2117,G1086,G1166,G1171,G1172,G1173,
     G1174,G1175,G1176,G1177,G1178,G1179,G1181,G1182,G1183,G1184,G1188,
     G1189,G1190,G1191,G1192,G1193,G1194,G1195,G1196,G1197,G1437,G1442,
     G1443,G1444,G1445,G1446,G1447,G1451,G1454,G1455,G1456,G1457,G1465,
     G1466,G1467,G1468,G1469,G1470,G1471,G1472,G1473,G1474,G1475,G1476,
     G1477,G1481,G1482,G1764,G1843,G1850,G1851,G1853,G1854,G1855,G1856,
     G1857,G1859,G1860,G1861,G1862,G1867,G1868,G1869,G1870,G1871,G1872,
     G1873,G1874,G1878,G2113,G2120,G2121,G2123,G2124,G2128,G2131,G2132,
     G2133,G2134,G2143,G2144,G2145,G2147,G2148,G2149,G2150,G2151,G2152,
     G2153,G2154,G2158,G2159,G3449,G3458,G3472,G3481,G3497,G3501,G3505,
     G3509,G3531,G5428,G3967,G4191,G4199,G4207,G4215,G4223,G4231,G4239,
     G4247,G4255,G4263,G4271,G4371,G4381,G4391,G4401,G4429,G4439,G4449,
     G4459,G4497,G4507,G4517,G4527,G4537,G4547,G4585,G4595,G4605,G4615,
     G4719,G4727,G4735,G4751,G4759,G4835,G4845,G4893,G4903,G4961,G4971,
     G4981,G5049,G5059,G5069,G5222,G5223,G5232,G5233,G5294,G5395,G589,
     G616,G619,G627,G1185,G1448,G1458,G1478,G1863,G4747,G2125,G2135,
     G2155,G4995,G5005,G3533,G3921,G3925,G3929,G3933,G3943,G3946,G3949,
     G3952,G3966,G4107,G4196,G4204,G4212,G4220,G4244,G4252,G4260,G4268,
     G4361,G4419,G4467,G4487,G4555,G4575,G4684,G4692,G4700,G4708,G4732,
     G4740,G4748,G4825,G4883,G4928,G4941,G5009,G5029,G5224,G5225,G5234,
     G5235,G5376,G5417,G576,G1198,G4195,G4203,G4211,G4219,G4227,G1217,
     G4235,G1221,G4243,G1224,G4251,G4259,G4267,G4275,G1453,G4405,G4463,
     G4541,G4551,G1895,G4723,G1899,G4731,G1902,G4739,G4755,G1929,G4763,
     G2130,G3500,G3504,G3508,G3512,G3520,G3523,G3526,G3529,G3837,G3942,
     G3945,G3948,G3951,G3968,G4375,G4385,G4395,G4433,G4443,G4453,G4501,
     G4511,G4521,G4531,G4619,G4589,G4599,G4609,G4839,G4849,G4897,G4907,
     G4965,G4975,G4985,G5073,G5053,G5063,G5247,G5255,G590,G617,G620,
     G628,G3535,G1199,G4202,G1204,G4210,G1207,G4218,G1211,G4226,G1214,
     G1218,G1222,G1225,G4250,G1237,G4258,G1242,G4266,G1247,G4274,G1252,
     G1462,G4690,G1882,G4698,G1885,G4706,G1889,G4714,G1892,G1896,G1900,
     G1903,G4738,G1915,G4746,G1920,G4754,G1925,G1930,G2139,G3519,G3522,
     G3525,G3528,G3848,G3944,G3947,G3950,G3953,G5421,G4111,G4112,G4351,
     G4365,G4409,G4423,G4471,G4472,G4477,G4491,G4559,G4560,G4565,G4579,
     G4815,G4829,G4873,G4887,G4931,G4934,G4945,G5013,G5014,G5019,G5033,
     G5382,G5385,G3970,G1200,G1203,G1206,G1210,G1213,G1219,G1223,G1236,
     G1241,G1246,G1251,G1881,G1884,G1888,G1891,G1897,G1901,G1914,G1919,
     G1924,G1931,G3521,G3524,G3527,G3530,G5251,G5259,G4113,G4473,G4561,
     G5015,G5384,G5406,G5414,G1664,G2335,G718,G855,G1205,G1208,G1212,
     G1215,G1220,G1231,G1238,G1243,G1248,G1253,G1272,G1483,G1883,G1886,
     G1890,G1893,G1898,G1909,G1916,G1921,G1926,G1953,G2160,G4355,G4356,
     G4413,G4414,G4474,G4481,G4562,G4569,G4819,G4820,G4877,G4878,G4935,
     G4936,G5016,G5023,G5244,G5252,G5409,G566,G577,G3733,G1209,G1216,
     G1257,G1262,G1267,G1887,G1894,G1935,G1943,G1948,G3779,G3840,G5412,
     G5420,G3964,G4357,G4415,G4821,G4879,G4937,G567,G568,G569,G570,
     G578,G579,G580,G1256,G1261,G1266,G1271,G1486,G1934,G1942,G1947,
     G1952,G2163,G5250,G3537,G5258,G3542,G3782,G3785,G3788,G3790,G3843,
     G3846,G3849,G3960,G5413,G3963,G4010,G4068,G4358,G4416,G4480,G4483,
     G4568,G4571,G4822,G4880,G4938,G5022,G5025,G1258,G1263,G1268,G1273,
     G1936,G1944,G1949,G1954,G3536,G3541,G3791,G3792,G3793,G3850,G3851,
     G3961,G3965,G4024,G4082,G4482,G4570,G5024,G1666,G1670,G2337,G2341,
     G719,G758,G798,G856,G3538,G3543,G3962,G4364,G4367,G4422,G4425,
     G4484,G4572,G4828,G4831,G4886,G4889,G4944,G4947,G5026,G571,G572,
     G573,G574,G581,G582,G583,G584,G1576,G1578,G659,G1672,G1676,
     G1678,G1682,G1684,G2250,G2252,G691,G2343,G2347,G2349,G2353,G2355,
     G743,G744,G748,G749,G753,G754,G759,G783,G784,G788,G789,
     G793,G794,G799,G3735,G3835,G3651,G4013,G4016,G4019,G4022,G4071,
     G4074,G4077,G4080,G4096,G4366,G4424,G4830,G4888,G4946,G640,G662,
     G665,G668,G674,G694,G697,G700,G817,G839,G3540,G3545,G3777,
     G3648,G4025,G4026,G4027,G4028,G4083,G4084,G4085,G4086,G4368,G4426,
     G4490,G4493,G4578,G4581,G4832,G4890,G4948,G5032,G5035,G811,G812,
     G853,G878,G4492,G4580,G5034,G1582,G1584,G1588,G1590,G1594,G1596,
     G1600,G1602,G2256,G2258,G2262,G2264,G2268,G2270,G2274,G2276,G708,
     G709,G723,G724,G728,G729,G733,G734,G738,G739,G768,G769,
     G773,G774,G778,G779,G4374,G4377,G4432,G4435,G4494,G4582,G4838,
     G4841,G4896,G4899,G4954,G4957,G5036,G643,G646,G649,G652,G677,
     G680,G683,G686,G4376,G4434,G4840,G4898,G4956,G4378,G4436,G4500,
     G4503,G4588,G4591,G4842,G4900,G4958,G5042,G5045,G4502,G4590,G5044,
     G4384,G4387,G4442,G4445,G4504,G4592,G4848,G4851,G4906,G4909,G4964,
     G4967,G5046,G4386,G4444,G4850,G4908,G4966,G4388,G4446,G4510,G4513,
     G4598,G4601,G4852,G4910,G4968,G5052,G5055,G4512,G4600,G5054,G4394,
     G4397,G4452,G4455,G4514,G4602,G4858,G4861,G4916,G4919,G4974,G4977,
     G5056,G4396,G4454,G4860,G4918,G4976,G4398,G4456,G4520,G4523,G4608,
     G4611,G4862,G4920,G4978,G5062,G5065,G4522,G4610,G5064,G4404,G1488,
     G4462,G1493,G4868,G2165,G4926,G2170,G4524,G4612,G4984,G4987,G5066,
     G1487,G1492,G2164,G2169,G4986,G1489,G1494,G2166,G2171,G4530,G4533,
     G4618,G4543,G4988,G5072,G4997,G4532,G4542,G4996,G1513,G1514,G1515,
     G1516,G4994,G2184,G2190,G2191,G2192,G2193,G4534,G4544,G4998,G2183,
     G4620,G5074,G4540,G1507,G4550,G1510,G2185,G5004,G2187,G1506,G1509,
     G4626,G2186,G2195,G5080,G1508,G1511,G2188,G1512,G1518,G2189,G1517,
     G2194,G4623,G5077,G1519,G4627,G2196,G5081,G1520,G2197,G1521,G2198,
     G840,G879,G1524,G2201,G3649,G3652,G3657,G3658,G3636,G3639,G3642,
     G3645,G3653,G3654,G3655,G3656,G763,G764,G803,G804,G1657,G1659,
     G2328,G2330,G1662,G2333,G657,G689,G1179_tmp,G1184_tmp,G1191_tmp,G1451_tmp,G1457_tmp,
     G1857_tmp,G1862_tmp,G1869_tmp,G2128_tmp,G2134_tmp,G1185_tmp,G1458_tmp,G1863_tmp,G2135_tmp,G4244_tmp,G4487_tmp,
     G4732_tmp,G4941_tmp,G575_0_tmp,G575_1_tmp,G585_0_tmp,G585_1_tmp,G853_tmp;

    buf g_G144 (G144, G141);
    buf g_G298 (G298, G293);
    and g_G4114 (G4114, G135, G4115);
    not g_G2825 (G2825, G2824);
    buf g_G973 (G973, G3173);
    not g_G3547 (G3547, G3546);
    not g_G3549 (G3549, G3548);
    not g_G3551 (G3551, G3550);
    not g_G3553 (G3553, G3552);
    not g_G594 (G594, G545);
    not g_G599 (G599, G348);
    not g_G600 (G600, G366);
    and g_G601 (G601, G552, G562);
    not g_G602 (G602, G549);
    not g_G603 (G603, G545);
    not g_G604 (G604, G545);
    not g_G611 (G611, G338);
    not g_G612 (G612, G358);
    nand g_G633 (G633, G373, G1);
    and g_G810 (G810, G141, G145);
    not g_G814 (G814, G3173);
    not g_G816 (G816, G4114);
    and g_G844 (G844, G2825, G27);
    and g_G846 (G846, G386, G556);
    not g_G848 (G848, G245);
    not g_G849 (G849, G552);
    not g_G850 (G850, G562);
    not g_G851 (G851, G559);
    and g_G852 (G852, G386, G559, G556, G552);
    not g_G1502 (G1502, G1497);
    buf g_G1528 (G1528, G1689);
    buf g_G1552 (G1552, G1690);
    buf g_G1609 (G1609, G1689);
    buf g_G1633 (G1633, G1690);
    buf g_G1697 (G1697, G137);
    buf g_G1698 (G1698, G137);
    buf g_G1701 (G1701, G141);
    not g_G2179 (G2179, G2174);
    buf g_G2203 (G2203, G1691);
    buf g_G2226 (G2226, G1694);
    buf g_G2281 (G2281, G1691);
    buf g_G2304 (G2304, G1694);
    buf g_G2361 (G2361, G254);
    buf g_G2370 (G2370, G251);
    buf g_G2382 (G2382, G251);
    buf g_G2393 (G2393, G248);
    buf g_G2405 (G2405, G248);
    buf g_G2418 (G2418, G4088);
    buf g_G2442 (G2442, G4087);
    buf g_G2476 (G2476, G4089);
    buf g_G2500 (G2500, G4090);
    buf g_G2533 (G2533, G210);
    buf g_G2537 (G2537, G210);
    buf g_G2541 (G2541, G218);
    buf g_G2545 (G2545, G218);
    buf g_G2549 (G2549, G226);
    buf g_G2553 (G2553, G226);
    buf g_G2557 (G2557, G234);
    buf g_G2561 (G2561, G234);
    buf g_G2627 (G2627, G257);
    buf g_G2631 (G2631, G257);
    buf g_G2635 (G2635, G265);
    buf g_G2639 (G2639, G265);
    buf g_G2643 (G2643, G273);
    buf g_G2647 (G2647, G273);
    buf g_G2651 (G2651, G281);
    buf g_G2655 (G2655, G281);
    buf g_G2721 (G2721, G335);
    buf g_G2734 (G2734, G335);
    buf g_G2816 (G2816, G206);
    and g_G2822 (G2822, G27, G31);
    buf g_G2826 (G2826, G1);
    buf g_G2828 (G2828, G2358);
    buf g_G2882 (G2882, G293);
    buf g_G2886 (G2886, G302);
    buf g_G2890 (G2890, G308);
    buf g_G2894 (G2894, G308);
    buf g_G2898 (G2898, G316);
    buf g_G2902 (G2902, G316);
    buf g_G2948 (G2948, G324);
    buf g_G2952 (G2952, G324);
    buf g_G2956 (G2956, G341);
    buf g_G2960 (G2960, G341);
    buf g_G2964 (G2964, G351);
    buf g_G2968 (G2968, G351);
    buf g_G3024 (G3024, G257);
    buf g_G3028 (G3028, G257);
    buf g_G3032 (G3032, G265);
    buf g_G3036 (G3036, G265);
    buf g_G3040 (G3040, G273);
    buf g_G3044 (G3044, G273);
    buf g_G3048 (G3048, G281);
    buf g_G3052 (G3052, G281);
    buf g_G3092 (G3092, G332);
    buf g_G3105 (G3105, G332);
    buf g_G3175 (G3175, G549);
    and g_G3176 (G3176, G31, G27);
    not g_G3181 (G3181, G2358);
    buf g_G3204 (G3204, G324);
    buf g_G3208 (G3208, G324);
    buf g_G3212 (G3212, G341);
    buf g_G3216 (G3216, G341);
    buf g_G3220 (G3220, G351);
    buf g_G3224 (G3224, G351);
    buf g_G3256 (G3256, G293);
    buf g_G3260 (G3260, G302);
    buf g_G3264 (G3264, G308);
    buf g_G3268 (G3268, G308);
    buf g_G3272 (G3272, G316);
    buf g_G3276 (G3276, G316);
    buf g_G3302 (G3302, G361);
    buf g_G3314 (G3314, G361);
    buf g_G3354 (G3354, G210);
    buf g_G3358 (G3358, G210);
    buf g_G3362 (G3362, G218);
    buf g_G3366 (G3366, G218);
    buf g_G3370 (G3370, G226);
    buf g_G3374 (G3374, G226);
    buf g_G3378 (G3378, G234);
    buf g_G3382 (G3382, G234);
    not g_G3440 (G3440, G324);
    buf g_G3554 (G3554, G242);
    buf g_G3555 (G3555, G242);
    buf g_G3556 (G3556, G254);
    buf g_G3558 (G3558, G4088);
    buf g_G3582 (G3582, G4087);
    buf g_G3616 (G3616, G4092);
    buf g_G3628 (G3628, G4091);
    buf g_G3660 (G3660, G4089);
    buf g_G3684 (G3684, G4090);
    not g_G3721 (G3721, G3717);
    not g_G3728 (G3728, G3724);
    buf g_G3737 (G3737, G4091);
    buf g_G3757 (G3757, G4092);
    buf g_G3795 (G3795, G4091);
    buf g_G3815 (G3815, G4092);
    buf g_G3972 (G3972, G4091);
    buf g_G3991 (G3991, G4092);
    buf g_G4030 (G4030, G4091);
    buf g_G4049 (G4049, G4092);
    buf g_G4110 (G4110, G299);
    buf g_G4119 (G4119, G446);
    buf g_G4127 (G4127, G457);
    buf g_G4135 (G4135, G468);
    buf g_G4143 (G4143, G422);
    buf g_G4151 (G4151, G435);
    buf g_G4159 (G4159, G389);
    buf g_G4167 (G4167, G400);
    buf g_G4175 (G4175, G411);
    buf g_G4183 (G4183, G374);
    buf g_G4188 (G4188, G4);
    buf g_G4276 (G4276, G446);
    buf g_G4284 (G4284, G457);
    buf g_G4292 (G4292, G468);
    buf g_G4300 (G4300, G435);
    buf g_G4308 (G4308, G389);
    buf g_G4316 (G4316, G400);
    buf g_G4324 (G4324, G411);
    buf g_G4332 (G4332, G422);
    buf g_G4340 (G4340, G374);
    buf g_G4631 (G4631, G479);
    buf g_G4639 (G4639, G490);
    buf g_G4647 (G4647, G503);
    buf g_G4655 (G4655, G514);
    buf g_G4663 (G4663, G523);
    buf g_G4671 (G4671, G534);
    buf g_G4676 (G4676, G54);
    buf g_G4764 (G4764, G479);
    buf g_G4772 (G4772, G503);
    buf g_G4780 (G4780, G514);
    buf g_G4788 (G4788, G523);
    buf g_G4796 (G4796, G534);
    buf g_G4804 (G4804, G490);
    buf g_G5082 (G5082, G361);
    buf g_G5085 (G5085, G369);
    buf g_G5090 (G5090, G341);
    buf g_G5093 (G5093, G351);
    buf g_G5098 (G5098, G308);
    buf g_G5101 (G5101, G316);
    buf g_G5108 (G5108, G293);
    buf g_G5111 (G5111, G302);
    buf g_G5332 (G5332, G281);
    buf g_G5335 (G5335, G289);
    buf g_G5340 (G5340, G265);
    buf g_G5343 (G5343, G273);
    buf g_G5348 (G5348, G234);
    buf g_G5351 (G5351, G257);
    buf g_G5356 (G5356, G218);
    buf g_G5359 (G5359, G226);
    buf g_G5369 (G5369, G210);
    not g_G634 (G634, G633);
    and g_G815 (G815, G136, G814);
    not g_G845 (G845, G844);
    not g_G847 (G847, G846);
    buf g_G926 (G926, G1697);
    buf g_G923 (G923, G1701);
    buf g_G921 (G921, G2826);
    and g_G2979 (G2979, G3553, G514);
    or g_G2999 (G2999, G3547, G514);
    buf g_G892 (G892, G3175);
    buf g_G887 (G887, G4110);
    not g_G606 (G606, G3175);
    and g_G1580 (G1580, G170, G1528, G1552);
    and g_G1586 (G1586, G173, G1528, G1552);
    and g_G1592 (G1592, G167, G1528, G1552);
    and g_G1598 (G1598, G164, G1528, G1552);
    and g_G1604 (G1604, G161, G1528, G1552);
    nand g_G656 (G656, G2822, G140);
    and g_G1668 (G1668, G185, G1609, G1633);
    and g_G1674 (G1674, G158, G1609, G1633);
    and g_G1680 (G1680, G152, G1609, G1633);
    and g_G1686 (G1686, G146, G1609, G1633);
    and g_G2254 (G2254, G170, G2203, G2226);
    and g_G2260 (G2260, G173, G2203, G2226);
    and g_G2266 (G2266, G167, G2203, G2226);
    and g_G2272 (G2272, G164, G2203, G2226);
    and g_G2278 (G2278, G161, G2203, G2226);
    and g_G2339 (G2339, G185, G2281, G2304);
    and g_G2345 (G2345, G158, G2281, G2304);
    and g_G2351 (G2351, G152, G2281, G2304);
    and g_G2357 (G2357, G146, G2281, G2304);
    and g_G711 (G711, G106, G3660, G3684);
    and g_G721 (G721, G61, G2418, G2442);
    and g_G726 (G726, G106, G3558, G3582);
    and g_G731 (G731, G49, G3558, G3582);
    and g_G736 (G736, G103, G3558, G3582);
    and g_G741 (G741, G40, G3558, G3582);
    and g_G746 (G746, G37, G3558, G3582);
    and g_G751 (G751, G20, G2418, G2442);
    and g_G756 (G756, G17, G2418, G2442);
    and g_G761 (G761, G70, G2418, G2442);
    and g_G766 (G766, G64, G2418, G2442);
    and g_G771 (G771, G49, G3660, G3684);
    and g_G776 (G776, G103, G3660, G3684);
    and g_G781 (G781, G40, G3660, G3684);
    and g_G786 (G786, G37, G3660, G3684);
    and g_G791 (G791, G20, G2476, G2500);
    and g_G796 (G796, G17, G2476, G2500);
    and g_G801 (G801, G70, G2476, G2500);
    and g_G806 (G806, G64, G2476, G2500);
    not g_G809 (G809, G2822);
    and g_G3734 (G3734, G123, G3728, G3717);
    and g_G842 (G842, G3795, G3815);
    and g_G858 (G858, G61, G2476, G2500);
    and g_G881 (G881, G3737, G3757);
    not g_G4123 (G4123, G4119);
    not g_G4131 (G4131, G4127);
    not g_G4139 (G4139, G4135);
    not g_G4147 (G4147, G4143);
    not g_G4155 (G4155, G4151);
    not g_G4163 (G4163, G4159);
    not g_G4171 (G4171, G4167);
    not g_G4179 (G4179, G4175);
    not g_G4187 (G4187, G4183);
    not g_G4194 (G4194, G4188);
    not g_G4282 (G4282, G4276);
    not g_G4290 (G4290, G4284);
    not g_G4298 (G4298, G4292);
    not g_G4306 (G4306, G4300);
    not g_G4314 (G4314, G4308);
    not g_G4322 (G4322, G4316);
    not g_G4330 (G4330, G4324);
    not g_G4338 (G4338, G4332);
    not g_G4346 (G4346, G4340);
    buf g_G1526 (G1526, G1697);
    not g_G1540 (G1540, G1528);
    not g_G1564 (G1564, G1552);
    buf g_G1606 (G1606, G1697);
    not g_G1621 (G1621, G1609);
    not g_G1645 (G1645, G1633);
    and g_G1661 (G1661, G179, G1609, G1633);
    buf g_G1688 (G1688, G2826);
    not g_G4635 (G4635, G4631);
    not g_G4643 (G4643, G4639);
    not g_G4651 (G4651, G4647);
    not g_G4659 (G4659, G4655);
    not g_G4667 (G4667, G4663);
    not g_G4675 (G4675, G4671);
    not g_G4682 (G4682, G4676);
    not g_G4770 (G4770, G4764);
    not g_G4778 (G4778, G4772);
    not g_G4786 (G4786, G4780);
    not g_G4794 (G4794, G4788);
    not g_G4802 (G4802, G4796);
    not g_G4810 (G4810, G4804);
    buf g_G2202 (G2202, G1698);
    not g_G2215 (G2215, G2203);
    not g_G2238 (G2238, G2226);
    buf g_G2279 (G2279, G1698);
    not g_G2293 (G2293, G2281);
    not g_G2316 (G2316, G2304);
    and g_G2332 (G2332, G179, G2281, G2304);
    not g_G2430 (G2430, G2418);
    not g_G2454 (G2454, G2442);
    not g_G2488 (G2488, G2476);
    not g_G2512 (G2512, G2500);
    not g_G2536 (G2536, G2533);
    not g_G2540 (G2540, G2537);
    not g_G2544 (G2544, G2541);
    not g_G2548 (G2548, G2545);
    not g_G2552 (G2552, G2549);
    not g_G2556 (G2556, G2553);
    not g_G2560 (G2560, G2557);
    not g_G2564 (G2564, G2561);
    and g_G2566 (G2566, G3553, G457, G2537);
    and g_G2572 (G2572, G3553, G468, G2545);
    and g_G2578 (G2578, G3553, G422, G2553);
    and g_G2584 (G2584, G3553, G435, G2561);
    and g_G2590 (G2590, G3547, G2533);
    and g_G2595 (G2595, G3547, G2541);
    and g_G2600 (G2600, G3547, G2549);
    and g_G2605 (G2605, G3547, G2557);
    not g_G2630 (G2630, G2627);
    not g_G2634 (G2634, G2631);
    not g_G2638 (G2638, G2635);
    not g_G2642 (G2642, G2639);
    not g_G2646 (G2646, G2643);
    not g_G2650 (G2650, G2647);
    not g_G2654 (G2654, G2651);
    not g_G2658 (G2658, G2655);
    and g_G2660 (G2660, G3553, G389, G2631);
    and g_G2666 (G2666, G3553, G400, G2639);
    and g_G2672 (G2672, G3553, G411, G2647);
    and g_G2678 (G2678, G3553, G374, G2655);
    and g_G2684 (G2684, G3547, G2627);
    and g_G2689 (G2689, G3547, G2635);
    and g_G2694 (G2694, G3547, G2643);
    and g_G2699 (G2699, G3547, G2651);
    not g_G2728 (G2728, G2721);
    not g_G2741 (G2741, G2734);
    and g_G2748 (G2748, G292, G2721);
    and g_G2750 (G2750, G288, G2721);
    and g_G2752 (G2752, G280, G2721);
    and g_G2754 (G2754, G272, G2721);
    and g_G2756 (G2756, G264, G2721);
    and g_G2758 (G2758, G241, G2734);
    and g_G2760 (G2760, G233, G2734);
    and g_G2762 (G2762, G225, G2734);
    and g_G2764 (G2764, G217, G2734);
    and g_G2766 (G2766, G209, G2734);
    buf g_G2827 (G2827, G1701);
    not g_G2838 (G2838, G2828);
    not g_G2847 (G2847, G2822);
    not g_G2885 (G2885, G2882);
    not g_G2889 (G2889, G2886);
    not g_G2893 (G2893, G2890);
    not g_G2897 (G2897, G2894);
    not g_G2901 (G2901, G2898);
    not g_G2905 (G2905, G2902);
    and g_G2906 (G2906, G2393, G2886);
    and g_G2909 (G2909, G2393, G479, G2894);
    and g_G2913 (G2913, G2393, G490, G2902);
    and g_G2918 (G2918, G3554, G2882);
    and g_G2922 (G2922, G3554, G2890);
    and g_G2927 (G2927, G3554, G2898);
    not g_G2951 (G2951, G2948);
    not g_G2955 (G2955, G2952);
    not g_G2959 (G2959, G2956);
    not g_G2963 (G2963, G2960);
    not g_G2967 (G2967, G2964);
    not g_G2971 (G2971, G2968);
    and g_G2973 (G2973, G3553, G503, G2952);
    not g_G2980 (G2980, G2979);
    and g_G2982 (G2982, G3553, G523, G2960);
    and g_G2988 (G2988, G3553, G534, G2968);
    and g_G2994 (G2994, G3547, G2948);
    and g_G3001 (G3001, G3547, G2956);
    and g_G3006 (G3006, G3547, G2964);
    not g_G3027 (G3027, G3024);
    not g_G3031 (G3031, G3028);
    not g_G3035 (G3035, G3032);
    not g_G3039 (G3039, G3036);
    not g_G3043 (G3043, G3040);
    not g_G3047 (G3047, G3044);
    not g_G3051 (G3051, G3048);
    not g_G3055 (G3055, G3052);
    and g_G3056 (G3056, G2393, G389, G3028);
    and g_G3060 (G3060, G2393, G400, G3036);
    and g_G3064 (G3064, G2393, G411, G3044);
    and g_G3068 (G3068, G2393, G374, G3052);
    and g_G3073 (G3073, G3554, G3024);
    and g_G3078 (G3078, G3554, G3032);
    and g_G3083 (G3083, G3554, G3040);
    and g_G3088 (G3088, G3554, G3048);
    not g_G3099 (G3099, G3092);
    not g_G3112 (G3112, G3105);
    and g_G3119 (G3119, G372, G3092);
    and g_G3121 (G3121, G366, G3092);
    and g_G3123 (G3123, G358, G3092);
    and g_G3125 (G3125, G348, G3092);
    and g_G3126 (G3126, G338, G3092);
    and g_G3128 (G3128, G331, G3105);
    and g_G3130 (G3130, G323, G3105);
    and g_G3132 (G3132, G315, G3105);
    and g_G3134 (G3134, G307, G3105);
    and g_G3136 (G3136, G299, G3105);
    not g_G3187 (G3187, G3181);
    and g_G3193 (G3193, G83, G3181);
    and g_G3196 (G3196, G86, G3181);
    and g_G3199 (G3199, G88, G3181);
    and g_G3202 (G3202, G88, G3181);
    not g_G3207 (G3207, G3204);
    not g_G3211 (G3211, G3208);
    not g_G3215 (G3215, G3212);
    not g_G3219 (G3219, G3216);
    not g_G3223 (G3223, G3220);
    not g_G3227 (G3227, G3224);
    and g_G3228 (G3228, G2405, G503, G3208);
    and g_G3232 (G3232, G2405, G514);
    and g_G3234 (G3234, G2405, G523, G3216);
    and g_G3238 (G3238, G2405, G534, G3224);
    and g_G3243 (G3243, G3555, G3204);
    or g_G3247 (G3247, G3555, G514);
    and g_G3249 (G3249, G3555, G3212);
    and g_G3253 (G3253, G3555, G3220);
    not g_G3259 (G3259, G3256);
    not g_G3263 (G3263, G3260);
    not g_G3267 (G3267, G3264);
    not g_G3271 (G3271, G3268);
    not g_G3275 (G3275, G3272);
    not g_G3279 (G3279, G3276);
    and g_G3280 (G3280, G2405, G3260);
    and g_G3283 (G3283, G2405, G479, G3268);
    and g_G3287 (G3287, G2405, G490, G3276);
    and g_G3292 (G3292, G3555, G3256);
    and g_G3295 (G3295, G3555, G3264);
    and g_G3299 (G3299, G3555, G3272);
    not g_G3305 (G3305, G3302);
    buf g_G3306 (G3306, G2816);
    buf g_G3310 (G3310, G2816);
    not g_G3317 (G3317, G3314);
    buf g_G3318 (G3318, G2816);
    buf g_G3322 (G3322, G2816);
    and g_G3326 (G3326, G2405, G3302);
    and g_G3333 (G3333, G2405, G3314);
    not g_G3357 (G3357, G3354);
    not g_G3361 (G3361, G3358);
    not g_G3365 (G3365, G3362);
    not g_G3369 (G3369, G3366);
    not g_G3373 (G3373, G3370);
    not g_G3377 (G3377, G3374);
    not g_G3381 (G3381, G3378);
    not g_G3385 (G3385, G3382);
    and g_G3386 (G3386, G2393, G457, G3358);
    and g_G3390 (G3390, G2393, G468, G3366);
    and g_G3394 (G3394, G2393, G422, G3374);
    and g_G3398 (G3398, G2393, G435, G3382);
    and g_G3403 (G3403, G3554, G3354);
    and g_G3408 (G3408, G3554, G3362);
    and g_G3413 (G3413, G3554, G3370);
    and g_G3418 (G3418, G3554, G3378);
    not g_G5088 (G5088, G5082);
    not g_G5089 (G5089, G5085);
    not g_G5096 (G5096, G5090);
    not g_G5097 (G5097, G5093);
    buf g_G3489 (G3489, G3440);
    buf g_G3493 (G3493, G3440);
    not g_G3570 (G3570, G3558);
    not g_G3594 (G3594, G3582);
    not g_G3622 (G3622, G3616);
    not g_G3632 (G3632, G3628);
    and g_G3637 (G3637, G97, G3616);
    and g_G3640 (G3640, G94, G3616);
    and g_G3643 (G3643, G97, G3616);
    and g_G3646 (G3646, G94, G3616);
    not g_G3672 (G3672, G3660);
    not g_G3696 (G3696, G3684);
    not g_G3745 (G3745, G3737);
    not g_G3765 (G3765, G3757);
    not g_G3803 (G3803, G3795);
    not g_G3823 (G3823, G3815);
    not g_G5338 (G5338, G5332);
    not g_G5339 (G5339, G5335);
    not g_G5346 (G5346, G5340);
    not g_G5347 (G5347, G5343);
    not g_G5354 (G5354, G5348);
    not g_G5355 (G5355, G5351);
    not g_G3979 (G3979, G3972);
    not g_G3998 (G3998, G3991);
    not g_G4037 (G4037, G4030);
    not g_G4056 (G4056, G4049);
    buf g_G4094 (G4094, G4110);
    not g_G5104 (G5104, G5098);
    not g_G5105 (G5105, G5101);
    not g_G5114 (G5114, G5108);
    not g_G5115 (G5115, G5111);
    not g_G5362 (G5362, G5356);
    not g_G5363 (G5363, G5359);
    buf g_G5366 (G5366, G2816);
    not g_G5373 (G5373, G5369);
    buf g_G993 (G993, G1688);
    buf g_G978 (G978, G1688);
    buf g_G949 (G949, G1688);
    buf g_G939 (G939, G1688);
    and g_G2568 (G2568, G457, G3551, G2540);
    and g_G2574 (G2574, G468, G3551, G2548);
    and g_G2580 (G2580, G422, G3551, G2556);
    and g_G2586 (G2586, G435, G3551, G2564);
    and g_G2592 (G2592, G3549, G2536);
    and g_G2597 (G2597, G3549, G2544);
    and g_G2602 (G2602, G3549, G2552);
    and g_G2607 (G2607, G3549, G2560);
    and g_G2662 (G2662, G389, G3551, G2634);
    and g_G2668 (G2668, G400, G3551, G2642);
    and g_G2674 (G2674, G411, G3551, G2650);
    and g_G2680 (G2680, G374, G3551, G2658);
    and g_G2686 (G2686, G3549, G2630);
    and g_G2691 (G2691, G3549, G2638);
    and g_G2696 (G2696, G3549, G2646);
    and g_G2701 (G2701, G3549, G2654);
    and g_G2907 (G2907, G2370, G2889);
    and g_G2910 (G2910, G479, G2370, G2897);
    and g_G2914 (G2914, G490, G2370, G2905);
    and g_G2920 (G2920, G3556, G2885);
    and g_G2924 (G2924, G3556, G2893);
    and g_G2929 (G2929, G3556, G2901);
    and g_G2975 (G2975, G503, G3551, G2955);
    and g_G2984 (G2984, G523, G3551, G2963);
    and g_G2990 (G2990, G534, G3551, G2971);
    and g_G2996 (G2996, G3549, G2951);
    and g_G3003 (G3003, G3549, G2959);
    and g_G3008 (G3008, G3549, G2967);
    and g_G3015 (G3015, G2980, G2999);
    and g_G3057 (G3057, G389, G2370, G3031);
    and g_G3061 (G3061, G400, G2370, G3039);
    and g_G3065 (G3065, G411, G2370, G3047);
    and g_G3069 (G3069, G374, G2370, G3055);
    and g_G3075 (G3075, G3556, G3027);
    and g_G3080 (G3080, G3556, G3035);
    and g_G3085 (G3085, G3556, G3043);
    and g_G3090 (G3090, G3556, G3051);
    and g_G3229 (G3229, G503, G2382, G3211);
    not g_G3233 (G3233, G3232);
    and g_G3235 (G3235, G523, G2382, G3219);
    and g_G3239 (G3239, G534, G2382, G3227);
    and g_G3244 (G3244, G2361, G3207);
    and g_G3250 (G3250, G2361, G3215);
    and g_G3254 (G3254, G2361, G3223);
    and g_G3281 (G3281, G2382, G3263);
    and g_G3284 (G3284, G479, G2382, G3271);
    and g_G3288 (G3288, G490, G2382, G3279);
    and g_G3293 (G3293, G2361, G3259);
    and g_G3296 (G3296, G2361, G3267);
    and g_G3300 (G3300, G2361, G3275);
    and g_G3327 (G3327, G2382, G3305);
    and g_G3334 (G3334, G2382, G3317);
    and g_G3387 (G3387, G457, G2370, G3361);
    and g_G3391 (G3391, G468, G2370, G3369);
    and g_G3395 (G3395, G422, G2370, G3377);
    and g_G3399 (G3399, G435, G2370, G3385);
    and g_G3405 (G3405, G3556, G3357);
    and g_G3410 (G3410, G3556, G3365);
    and g_G3415 (G3415, G3556, G3373);
    and g_G3420 (G3420, G3556, G3381);
    nand g_G3422 (G3422, G5085, G5088);
    nand g_G3423 (G3423, G5082, G5089);
    nand g_G3431 (G3431, G5093, G5096);
    nand g_G3432 (G3432, G5090, G5097);
    nand g_G3895 (G3895, G5335, G5338);
    nand g_G3896 (G3896, G5332, G5339);
    nand g_G3904 (G3904, G5343, G5346);
    nand g_G3905 (G3905, G5340, G5347);
    nand g_G3913 (G3913, G5351, G5354);
    nand g_G3914 (G3914, G5348, G5355);
    buf g_G889 (G889, G4094);
    nand g_G5106 (G5106, G5101, G5104);
    nand g_G5107 (G5107, G5098, G5105);
    nand g_G5116 (G5116, G5111, G5114);
    nand g_G5117 (G5117, G5108, G5115);
    nand g_G5364 (G5364, G5359, G5362);
    nand g_G5365 (G5365, G5356, G5363);
    not g_G593 (G593, G4094);
    and g_G2880 (G2880, G2838, G2847);
    and g_G2881 (G2881, G2828, G2847);
    and g_G1579 (G1579, G200, G1540, G1552);
    and g_G1585 (G1585, G203, G1540, G1552);
    and g_G1591 (G1591, G197, G1540, G1552);
    and g_G1597 (G1597, G194, G1540, G1552);
    and g_G1603 (G1603, G191, G1540, G1552);
    and g_G1667 (G1667, G182, G1621, G1633);
    and g_G1673 (G1673, G188, G1621, G1633);
    and g_G1679 (G1679, G155, G1621, G1633);
    and g_G1685 (G1685, G149, G1621, G1633);
    and g_G2876 (G2876, G2838, G2847);
    and g_G2877 (G2877, G2828, G2847);
    and g_G2253 (G2253, G200, G2215, G2226);
    and g_G2259 (G2259, G203, G2215, G2226);
    and g_G2265 (G2265, G197, G2215, G2226);
    and g_G2271 (G2271, G194, G2215, G2226);
    and g_G2277 (G2277, G191, G2215, G2226);
    and g_G2338 (G2338, G182, G2293, G2304);
    and g_G2344 (G2344, G188, G2293, G2304);
    and g_G2350 (G2350, G155, G2293, G2304);
    and g_G2356 (G2356, G149, G2293, G2304);
    and g_G2868 (G2868, G2838, G2847);
    and g_G2869 (G2869, G2828, G2847);
    and g_G710 (G710, G109, G3672, G3684);
    and g_G2872 (G2872, G2838, G2847);
    and g_G2873 (G2873, G2828, G2847);
    and g_G720 (G720, G11, G2430, G2442);
    and g_G725 (G725, G109, G3570, G3582);
    and g_G730 (G730, G46, G3570, G3582);
    and g_G735 (G735, G100, G3570, G3582);
    and g_G740 (G740, G91, G3570, G3582);
    and g_G745 (G745, G43, G3570, G3582);
    and g_G750 (G750, G76, G2430, G2442);
    and g_G755 (G755, G73, G2430, G2442);
    and g_G760 (G760, G67, G2430, G2442);
    and g_G765 (G765, G14, G2430, G2442);
    and g_G770 (G770, G46, G3672, G3684);
    and g_G775 (G775, G100, G3672, G3684);
    and g_G780 (G780, G91, G3672, G3684);
    and g_G785 (G785, G43, G3672, G3684);
    and g_G790 (G790, G76, G2488, G2500);
    and g_G795 (G795, G73, G2488, G2500);
    and g_G800 (G800, G67, G2488, G2500);
    and g_G805 (G805, G14, G2488, G2500);
    and g_G841 (G841, G120, G3803, G3815);
    and g_G857 (G857, G11, G2488, G2500);
    and g_G880 (G880, G118, G3745, G3757);
    and g_G1660 (G1660, G176, G1621, G1633);
    and g_G2331 (G2331, G176, G2293, G2304);
    or g_G2569 (G2569, G2566, G2568);
    or g_G2575 (G2575, G2572, G2574);
    or g_G2581 (G2581, G2578, G2580);
    or g_G2587 (G2587, G2584, G2586);
    or g_G2593 (G2593, G2590, G2592, G457);
    or g_G2598 (G2598, G2595, G2597, G468);
    or g_G2603 (G2603, G2600, G2602, G422);
    or g_G2608 (G2608, G2605, G2607, G435);
    or g_G2663 (G2663, G2660, G2662);
    or g_G2669 (G2669, G2666, G2668);
    or g_G2675 (G2675, G2672, G2674);
    or g_G2681 (G2681, G2678, G2680);
    or g_G2687 (G2687, G2684, G2686, G389);
    or g_G2692 (G2692, G2689, G2691, G400);
    or g_G2697 (G2697, G2694, G2696, G411);
    or g_G2702 (G2702, G2699, G2701, G374);
    and g_G2747 (G2747, G289, G2728);
    and g_G2749 (G2749, G281, G2728);
    and g_G2751 (G2751, G273, G2728);
    and g_G2753 (G2753, G265, G2728);
    and g_G2755 (G2755, G257, G2728);
    and g_G2757 (G2757, G234, G2741);
    and g_G2759 (G2759, G226, G2741);
    and g_G2761 (G2761, G218, G2741);
    and g_G2763 (G2763, G210, G2741);
    and g_G2765 (G2765, G206, G2741);
    not g_G2857 (G2857, G2847);
    or g_G2908 (G2908, G2906, G2907);
    or g_G2911 (G2911, G2909, G2910);
    or g_G2915 (G2915, G2913, G2914);
    or g_G2925 (G2925, G2922, G2924, G479);
    or g_G2930 (G2930, G2927, G2929, G490);
    or g_G2933 (G2933, G2918, G2920);
    or g_G2976 (G2976, G2973, G2975);
    or g_G2985 (G2985, G2982, G2984);
    or g_G2991 (G2991, G2988, G2990);
    or g_G2997 (G2997, G2994, G2996, G503);
    or g_G3004 (G3004, G3001, G3003, G523);
    or g_G3009 (G3009, G3006, G3008, G534);
    or g_G3058 (G3058, G3056, G3057);
    or g_G3062 (G3062, G3060, G3061);
    or g_G3066 (G3066, G3064, G3065);
    or g_G3070 (G3070, G3068, G3069);
    or g_G3076 (G3076, G3073, G3075, G389);
    or g_G3081 (G3081, G3078, G3080, G400);
    or g_G3086 (G3086, G3083, G3085, G411);
    or g_G3091 (G3091, G3088, G3090, G374);
    and g_G3118 (G3118, G369, G3099);
    and g_G3120 (G3120, G361, G3099);
    and g_G3122 (G3122, G351, G3099);
    and g_G3124 (G3124, G341, G3099);
    and g_G3127 (G3127, G324, G3112);
    and g_G3129 (G3129, G316, G3112);
    and g_G3131 (G3131, G308, G3112);
    and g_G3133 (G3133, G302, G3112);
    and g_G3135 (G3135, G293, G3112);
    or g_G3147 (G3147, G3099, G3126);
    and g_G3192 (G3192, G83, G3187);
    and g_G3195 (G3195, G87, G3187);
    and g_G3198 (G3198, G34, G3187);
    and g_G3201 (G3201, G34, G3187);
    or g_G3230 (G3230, G3228, G3229);
    or g_G3236 (G3236, G3234, G3235);
    or g_G3240 (G3240, G3238, G3239);
    or g_G3245 (G3245, G3243, G3244, G503);
    or g_G3251 (G3251, G3249, G3250, G523);
    or g_G3255 (G3255, G3253, G3254, G534);
    or g_G3282 (G3282, G3280, G3281);
    or g_G3285 (G3285, G3283, G3284);
    or g_G3289 (G3289, G3287, G3288);
    or g_G3297 (G3297, G3295, G3296, G479);
    or g_G3301 (G3301, G3299, G3300, G490);
    not g_G3309 (G3309, G3306);
    not g_G3313 (G3313, G3310);
    not g_G3321 (G3321, G3318);
    not g_G3325 (G3325, G3322);
    or g_G3328 (G3328, G3326, G3327);
    and g_G3329 (G3329, G2405, G446, G3310);
    or g_G3335 (G3335, G3333, G3334);
    and g_G3336 (G3336, G2405, G446, G3322);
    and g_G3341 (G3341, G3555, G3306);
    and g_G3345 (G3345, G3555, G3318);
    or g_G3388 (G3388, G3386, G3387);
    or g_G3392 (G3392, G3390, G3391);
    or g_G3396 (G3396, G3394, G3395);
    or g_G3400 (G3400, G3398, G3399);
    or g_G3406 (G3406, G3403, G3405, G457);
    or g_G3411 (G3411, G3408, G3410, G468);
    or g_G3416 (G3416, G3413, G3415, G422);
    or g_G3421 (G3421, G3418, G3420, G435);
    nand g_G3424 (G3424, G3422, G3423);
    nand g_G3433 (G3433, G3431, G3432);
    not g_G3492 (G3492, G3489);
    not g_G3496 (G3496, G3493);
    and g_G3780 (G3780, G117, G3745, G3757);
    and g_G3783 (G3783, G126, G3745, G3757);
    and g_G3786 (G3786, G127, G3745, G3757);
    and g_G3789 (G3789, G128, G3745, G3757);
    and g_G3838 (G3838, G131, G3803, G3815);
    and g_G3841 (G3841, G129, G3803, G3815);
    and g_G3844 (G3844, G119, G3803, G3815);
    and g_G3847 (G3847, G130, G3803, G3815);
    nand g_G3897 (G3897, G3895, G3896);
    nand g_G3906 (G3906, G3904, G3905);
    nand g_G3915 (G3915, G3913, G3914);
    and g_G4011 (G4011, G122, G3979, G3991);
    and g_G4014 (G4014, G113, G3979, G3991);
    and g_G4017 (G4017, G53, G3979, G3991);
    and g_G4020 (G4020, G114, G3979, G3991);
    and g_G4023 (G4023, G115, G3979, G3991);
    and g_G4069 (G4069, G52, G4037, G4049);
    and g_G4072 (G4072, G112, G4037, G4049);
    and g_G4075 (G4075, G116, G4037, G4049);
    and g_G4078 (G4078, G121, G4037, G4049);
    and g_G4081 (G4081, G123, G4037, G4049);
    nand g_G5206 (G5206, G5116, G5117);
    nand g_G5209 (G5209, G5106, G5107);
    and g_G5307 (G5307, G3233, G3247);
    or g_G5322 (G5322, G3292, G3293);
    not g_G5372 (G5372, G5366);
    nand g_G5375 (G5375, G5366, G5373);
    nand g_G5399 (G5399, G5364, G5365);
    not g_G2813 (G2813, G3015);
    or g_G3197 (G3197, G3195, G3196);
    or g_G3200 (G3200, G3198, G3199);
    or g_G3203 (G3203, G3201, G3202);
    or g_G3194 (G3194, G3192, G3193);
    not g_G2570 (G2570, G2569);
    not g_G2576 (G2576, G2575);
    not g_G2582 (G2582, G2581);
    not g_G2588 (G2588, G2587);
    not g_G2664 (G2664, G2663);
    not g_G2670 (G2670, G2669);
    not g_G2676 (G2676, G2675);
    not g_G2682 (G2682, G2681);
    or g_G2767 (G2767, G2749, G2750);
    or g_G2772 (G2772, G2751, G2752);
    or g_G2776 (G2776, G2753, G2754);
    or g_G2780 (G2780, G2755, G2756);
    or g_G2784 (G2784, G2757, G2758);
    or g_G2788 (G2788, G2759, G2760);
    or g_G2794 (G2794, G2761, G2762);
    or g_G2798 (G2798, G2763, G2764);
    or g_G2802 (G2802, G2765, G2766);
    not g_G2912 (G2912, G2911);
    not g_G2916 (G2916, G2915);
    not g_G2936 (G2936, G2908);
    not g_G2977 (G2977, G2976);
    not g_G2986 (G2986, G2985);
    not g_G2992 (G2992, G2991);
    not g_G3059 (G3059, G3058);
    not g_G3063 (G3063, G3062);
    not g_G3067 (G3067, G3066);
    not g_G3071 (G3071, G3070);
    or g_G3137 (G3137, G3120, G3121);
    or g_G3139 (G3139, G3122, G3123);
    or g_G3143 (G3143, G3124, G3125);
    or g_G3151 (G3151, G3127, G3128);
    or g_G3155 (G3155, G3129, G3130);
    or g_G3161 (G3161, G3131, G3132);
    or g_G3165 (G3165, G3133, G3134);
    or g_G3167 (G3167, G3135, G3136);
    not g_G3231 (G3231, G3230);
    not g_G3237 (G3237, G3236);
    not g_G3241 (G3241, G3240);
    not g_G3286 (G3286, G3285);
    not g_G3290 (G3290, G3289);
    and g_G3330 (G3330, G446, G2382, G3313);
    and g_G3337 (G3337, G446, G2382, G3325);
    and g_G3342 (G3342, G2361, G3309);
    and g_G3346 (G3346, G2361, G3321);
    not g_G3348 (G3348, G3328);
    not g_G3352 (G3352, G3335);
    not g_G3389 (G3389, G3388);
    not g_G3393 (G3393, G3392);
    not g_G3397 (G3397, G3396);
    not g_G3401 (G3401, G3400);
    and g_G3845 (G3845, G3015, G3803, G3823);
    or g_G5126 (G5126, G3118, G3119);
    or g_G5178 (G5178, G2747, G2748);
    not g_G5325 (G5325, G3282);
    nand g_G5374 (G5374, G5369, G5372);
    not g_G2810 (G2810, G2933);
    and g_G635 (G635, G3197, G3176);
    and g_G2878 (G2878, G24, G2838, G2857);
    and g_G2879 (G2879, G25, G2828, G2857);
    and g_G2874 (G2874, G26, G2838, G2857);
    and g_G2875 (G2875, G81, G2828, G2857);
    and g_G703 (G703, G3200, G3176);
    and g_G2866 (G2866, G79, G2838, G2857);
    and g_G2867 (G2867, G23, G2828, G2857);
    and g_G2870 (G2870, G82, G2838, G2857);
    and g_G2871 (G2871, G80, G2828, G2857);
    and g_G716 (G716, G3203, G3176);
    and g_G819 (G819, G3194, G3176);
    and g_G1789 (G1789, G3147, G514);
    and g_G2036 (G2036, G514, G3147);
    and g_G2611 (G2611, G2570, G2593);
    and g_G2615 (G2615, G2576, G2598);
    and g_G2619 (G2619, G2582, G2603);
    and g_G2623 (G2623, G2588, G2608);
    and g_G2705 (G2705, G2664, G2687);
    and g_G2709 (G2709, G2670, G2692);
    and g_G2713 (G2713, G2676, G2697);
    and g_G2717 (G2717, G2682, G2702);
    and g_G2939 (G2939, G2912, G2925);
    and g_G2942 (G2942, G2916, G2930);
    buf g_G2945 (G2945, G2933);
    and g_G3012 (G3012, G2977, G2997);
    and g_G3018 (G3018, G2986, G3004);
    and g_G3021 (G3021, G2992, G3009);
    or g_G3331 (G3331, G3329, G3330);
    or g_G3338 (G3338, G3336, G3337);
    or g_G3343 (G3343, G3341, G3342, G446);
    or g_G3347 (G3347, G3345, G3346, G446);
    not g_G3428 (G3428, G3424);
    not g_G3437 (G3437, G3433);
    and g_G3514 (G3514, G3433, G3424, G3489);
    and g_G3836 (G3836, G3352, G3803, G3823);
    and g_G3852 (G3852, G3071, G3091);
    not g_G5311 (G5311, G5307);
    not g_G3901 (G3901, G3897);
    not g_G3910 (G3910, G3906);
    buf g_G3934 (G3934, G3915);
    buf g_G3938 (G3938, G3915);
    buf g_G4652 (G4652, G3147);
    buf g_G4783 (G4783, G3147);
    buf g_G5137 (G5137, G3147);
    not g_G5212 (G5212, G5206);
    not g_G5213 (G5213, G5209);
    and g_G5260 (G5260, G3063, G3081);
    and g_G5263 (G5263, G3067, G3086);
    and g_G5268 (G5268, G3401, G3421);
    and g_G5271 (G5271, G3059, G3076);
    and g_G5276 (G5276, G3393, G3411);
    and g_G5279 (G5279, G3397, G3416);
    and g_G5289 (G5289, G3389, G3406);
    and g_G5296 (G5296, G3237, G3251);
    and g_G5299 (G5299, G3241, G3255);
    and g_G5304 (G5304, G3231, G3245);
    and g_G5312 (G5312, G3286, G3297);
    and g_G5315 (G5315, G3290, G3301);
    not g_G5328 (G5328, G5322);
    nand g_G5396 (G5396, G5374, G5375);
    not g_G5403 (G5403, G5399);
    and g_G1286 (G1286, G446, G2802);
    not g_G2809 (G2809, G2936);
    not g_G597 (G597, G3348);
    and g_G1031 (G1031, G2802, G446);
    not g_G636 (G636, G635);
    or g_G637 (G637, G2878, G2879, G2880, G2881);
    or g_G671 (G671, G2874, G2875, G2876, G2877);
    not g_G704 (G704, G703);
    or g_G705 (G705, G2866, G2867, G2868, G2869);
    or g_G713 (G713, G2870, G2871, G2872, G2873);
    not g_G717 (G717, G716);
    not g_G820 (G820, G819);
    and g_G1046 (G1046, G2798, G457);
    and g_G1064 (G1064, G2794, G468);
    and g_G1071 (G1071, G422, G2788);
    and g_G1097 (G1097, G2784, G435);
    and g_G1111 (G1111, G2780, G389);
    and g_G1128 (G1128, G2776, G400);
    and g_G1145 (G1145, G2772, G411);
    and g_G1160 (G1160, G2767, G374);
    and g_G1301 (G1301, G457, G2798);
    and g_G1318 (G1318, G468, G2794);
    and g_G1324 (G1324, G422, G2788);
    and g_G1341 (G1341, G435, G2784);
    and g_G1359 (G1359, G389, G2780);
    and g_G1382 (G1382, G400, G2776);
    and g_G1404 (G1404, G411, G2772);
    and g_G1412 (G1412, G374, G2767);
    not g_G1704 (G1704, G3167);
    not g_G1712 (G1712, G3165);
    buf g_G1724 (G1724, G3165);
    and g_G1742 (G1742, G3161, G479);
    and g_G1749 (G1749, G490, G3155);
    and g_G1775 (G1775, G3151, G503);
    and g_G1806 (G1806, G3143, G523);
    and g_G1823 (G1823, G3139, G534);
    not g_G1829 (G1829, G3137);
    buf g_G1837 (G1837, G3137);
    not g_G1958 (G1958, G3167);
    not g_G1966 (G1966, G3165);
    buf g_G1978 (G1978, G3165);
    and g_G1995 (G1995, G479, G3161);
    and g_G2001 (G2001, G490, G3155);
    and g_G2018 (G2018, G503, G3151);
    and g_G2059 (G2059, G523, G3143);
    and g_G2081 (G2081, G534, G3139);
    buf g_G2089 (G2089, G3137);
    not g_G2106 (G2106, G3137);
    buf g_G3170 (G3170, G3167);
    not g_G3332 (G3332, G3331);
    not g_G3339 (G3339, G3338);
    not g_G5132 (G5132, G5126);
    not g_G5184 (G5184, G5178);
    not g_G3853 (G3853, G3852);
    not g_G3874 (G3874, G3348);
    and g_G4076 (G4076, G2936, G4037, G4056);
    buf g_G4116 (G4116, G2802);
    buf g_G4124 (G4124, G2798);
    buf g_G4132 (G4132, G2794);
    buf g_G4140 (G4140, G2788);
    buf g_G4148 (G4148, G2784);
    buf g_G4156 (G4156, G2780);
    buf g_G4164 (G4164, G2776);
    buf g_G4172 (G4172, G2772);
    buf g_G4180 (G4180, G2767);
    nor g_G4228 (G4228, G422, G2788);
    buf g_G4279 (G4279, G2802);
    buf g_G4287 (G4287, G2798);
    buf g_G4295 (G4295, G2794);
    buf g_G4303 (G4303, G2784);
    buf g_G4311 (G4311, G2780);
    buf g_G4319 (G4319, G2776);
    buf g_G4327 (G4327, G2772);
    buf g_G4335 (G4335, G2788);
    buf g_G4343 (G4343, G2767);
    nor g_G4348 (G4348, G422, G2788);
    nor g_G4464 (G4464, G374, G2767);
    buf g_G4628 (G4628, G3161);
    buf g_G4636 (G4636, G3155);
    buf g_G4644 (G4644, G3151);
    buf g_G4660 (G4660, G3143);
    buf g_G4668 (G4668, G3139);
    nor g_G4716 (G4716, G490, G3155);
    buf g_G4767 (G4767, G3161);
    buf g_G4775 (G4775, G3151);
    buf g_G4791 (G4791, G3143);
    buf g_G4799 (G4799, G3139);
    buf g_G4807 (G4807, G3155);
    nor g_G4812 (G4812, G490, G3155);
    buf g_G5118 (G5118, G3139);
    buf g_G5121 (G5121, G3143);
    buf g_G5129 (G5129, G3137);
    buf g_G5134 (G5134, G3151);
    buf g_G5142 (G5142, G3161);
    buf g_G5145 (G5145, G3155);
    buf g_G5152 (G5152, G3167);
    buf g_G5155 (G5155, G3165);
    buf g_G5162 (G5162, G2788);
    buf g_G5165 (G5165, G2784);
    buf g_G5170 (G5170, G2798);
    buf g_G5173 (G5173, G2794);
    buf g_G5181 (G5181, G2802);
    buf g_G5186 (G5186, G2772);
    buf g_G5189 (G5189, G2767);
    buf g_G5196 (G5196, G2780);
    buf g_G5199 (G5199, G2776);
    nand g_G5214 (G5214, G5209, G5212);
    nand g_G5215 (G5215, G5206, G5213);
    not g_G5329 (G5329, G5325);
    nand g_G5330 (G5330, G5325, G5328);
    not g_G2807 (G2807, G2942);
    not g_G2808 (G2808, G2939);
    not g_G2811 (G2811, G3021);
    not g_G2812 (G2812, G3018);
    not g_G2814 (G2814, G3012);
    not g_G2626 (G2626, G2623);
    not g_G2622 (G2622, G2619);
    not g_G2618 (G2618, G2615);
    not g_G2614 (G2614, G2611);
    not g_G2720 (G2720, G2717);
    not g_G2716 (G2716, G2713);
    not g_G2712 (G2712, G2709);
    not g_G2708 (G2708, G2705);
    and g_G639 (G639, G637, G2827);
    and g_G673 (G673, G671, G2827);
    and g_G707 (G707, G705, G2827);
    and g_G715 (G715, G713, G2827);
    and g_G3731 (G3731, G2945, G3728, G3721);
    not g_G4658 (G4658, G4652);
    nand g_G1777 (G1777, G4652, G4659);
    nand g_G2019 (G2019, G4783, G4786);
    not g_G4787 (G4787, G4783);
    and g_G3350 (G3350, G3332, G3343);
    and g_G3353 (G3353, G3339, G3347);
    not g_G5141 (G5141, G5137);
    and g_G3513 (G3513, G3428, G3433, G3492);
    and g_G3516 (G3516, G3424, G3437, G3496);
    and g_G3517 (G3517, G3437, G3428, G3493);
    and g_G3778 (G3778, G2717, G3745, G3765);
    and g_G3781 (G3781, G2713, G3745, G3765);
    and g_G3784 (G3784, G2709, G3745, G3765);
    and g_G3787 (G3787, G2705, G3745, G3765);
    and g_G3839 (G3839, G3021, G3803, G3823);
    and g_G3842 (G3842, G3018, G3803, G3823);
    not g_G5266 (G5266, G5260);
    not g_G5267 (G5267, G5263);
    not g_G5274 (G5274, G5268);
    not g_G5275 (G5275, G5271);
    not g_G5302 (G5302, G5296);
    not g_G5303 (G5303, G5299);
    not g_G5310 (G5310, G5304);
    nand g_G3891 (G3891, G5304, G5311);
    not g_G3937 (G3937, G3934);
    not g_G3941 (G3941, G3938);
    and g_G3955 (G3955, G3906, G3897, G3934);
    and g_G3958 (G3958, G3910, G3901, G3938);
    and g_G4009 (G4009, G2623, G3979, G3998);
    and g_G4012 (G4012, G2619, G3979, G3998);
    and g_G4015 (G4015, G2615, G3979, G3998);
    and g_G4018 (G4018, G2611, G3979, G3998);
    and g_G4067 (G4067, G3012, G4037, G4056);
    and g_G4070 (G4070, G2942, G4037, G4056);
    and g_G4073 (G4073, G2939, G4037, G4056);
    and g_G4079 (G4079, G2945, G4037, G4056);
    nand g_G5239 (G5239, G5214, G5215);
    not g_G5282 (G5282, G5276);
    not g_G5283 (G5283, G5279);
    not g_G5293 (G5293, G5289);
    not g_G5318 (G5318, G5312);
    not g_G5319 (G5319, G5315);
    nand g_G5331 (G5331, G5322, G5329);
    not g_G5402 (G5402, G5396);
    nand g_G5405 (G5405, G5396, G5403);
    and g_G595 (G595, G2807, G2808, G2809, G2810);
    and g_G596 (G596, G2811, G2812, G2813, G2814);
    and g_G607 (G607, G2626, G2622, G2618, G2614);
    and g_G608 (G608, G2720, G2716, G2712, G2708);
    and g_G1845 (G1845, G1704, G1724);
    and g_G1846 (G1846, G1712, G1704, G1742);
    and g_G2115 (G2115, G1958, G1978);
    and g_G2116 (G2116, G1966, G1958, G1995);
    not g_G4122 (G4122, G4116);
    nand g_G1022 (G1022, G4116, G4123);
    not g_G4130 (G4130, G4124);
    nand g_G1033 (G1033, G4124, G4131);
    not g_G4138 (G4138, G4132);
    nand g_G1051 (G1051, G4132, G4139);
    not g_G4146 (G4146, G4140);
    nand g_G1079 (G1079, G4140, G4147);
    not g_G4154 (G4154, G4148);
    nand g_G1088 (G1088, G4148, G4155);
    not g_G4162 (G4162, G4156);
    nand g_G1099 (G1099, G4156, G4163);
    not g_G4170 (G4170, G4164);
    nand g_G1115 (G1115, G4164, G4171);
    not g_G4178 (G4178, G4172);
    nand g_G1133 (G1133, G4172, G4179);
    not g_G4186 (G4186, G4180);
    nand g_G1151 (G1151, G4180, G4187);
    not g_G4234 (G4234, G4228);
    nand g_G1276 (G1276, G4279, G4282);
    not g_G4283 (G4283, G4279);
    nand g_G1287 (G1287, G4287, G4290);
    not g_G4291 (G4291, G4287);
    nand g_G1305 (G1305, G4295, G4298);
    not g_G4299 (G4299, G4295);
    nand g_G1330 (G1330, G4303, G4306);
    not g_G4307 (G4307, G4303);
    nand g_G1342 (G1342, G4311, G4314);
    not g_G4315 (G4315, G4311);
    nand g_G1363 (G1363, G4319, G4322);
    not g_G4323 (G4323, G4319);
    nand g_G1388 (G1388, G4327, G4330);
    not g_G4331 (G4331, G4327);
    nand g_G1420 (G1420, G4335, G4338);
    not g_G4339 (G4339, G4335);
    nand g_G1428 (G1428, G4343, G4346);
    not g_G4347 (G4347, G4343);
    not g_G4634 (G4634, G4628);
    nand g_G1729 (G1729, G4628, G4635);
    not g_G4642 (G4642, G4636);
    nand g_G1757 (G1757, G4636, G4643);
    not g_G4650 (G4650, G4644);
    nand g_G1766 (G1766, G4644, G4651);
    nand g_G1776 (G1776, G4655, G4658);
    not g_G4666 (G4666, G4660);
    nand g_G1793 (G1793, G4660, G4667);
    not g_G4674 (G4674, G4668);
    nand g_G1811 (G1811, G4668, G4675);
    and g_G1849 (G1849, G1712, G1742);
    and g_G1852 (G1852, G1712, G1742);
    and g_G1875 (G1875, G54, G1829);
    not g_G4722 (G4722, G4716);
    nand g_G1982 (G1982, G4767, G4770);
    not g_G4771 (G4771, G4767);
    nand g_G2007 (G2007, G4775, G4778);
    not g_G4779 (G4779, G4775);
    nand g_G2020 (G2020, G4780, G4787);
    nand g_G2040 (G2040, G4791, G4794);
    not g_G4795 (G4795, G4791);
    nand g_G2065 (G2065, G4799, G4802);
    not g_G4803 (G4803, G4799);
    nand g_G2097 (G2097, G4807, G4810);
    not g_G4811 (G4811, G4807);
    and g_G2119 (G2119, G1966, G1995);
    and g_G2122 (G2122, G1966, G1995);
    not g_G5124 (G5124, G5118);
    not g_G5125 (G5125, G5121);
    nand g_G3452 (G3452, G5129, G5132);
    not g_G5133 (G5133, G5129);
    not g_G5140 (G5140, G5134);
    nand g_G3462 (G3462, G5134, G5141);
    not g_G5168 (G5168, G5162);
    not g_G5169 (G5169, G5165);
    not g_G5176 (G5176, G5170);
    not g_G5177 (G5177, G5173);
    nand g_G3484 (G3484, G5181, G5184);
    not g_G5185 (G5185, G5181);
    nor g_G3515 (G3515, G3513, G3514);
    nor g_G3518 (G3518, G3516, G3517);
    not g_G3857 (G3857, G3853);
    nand g_G3860 (G3860, G5263, G5266);
    nand g_G3861 (G3861, G5260, G5267);
    nand g_G3869 (G3869, G5271, G5274);
    nand g_G3870 (G3870, G5268, G5275);
    not g_G3878 (G3878, G3874);
    nand g_G3881 (G3881, G5299, G5302);
    nand g_G3882 (G3882, G5296, G5303);
    nand g_G3890 (G3890, G5307, G5310);
    and g_G3954 (G3954, G3901, G3906, G3937);
    and g_G3957 (G3957, G3897, G3910, G3941);
    and g_G4021 (G4021, G3353, G3979, G3998);
    not g_G4099 (G4099, G3170);
    buf g_G4236 (G4236, G1071);
    not g_G4354 (G4354, G4348);
    buf g_G4406 (G4406, G1324);
    not g_G4470 (G4470, G4464);
    buf g_G4552 (G4552, G1412);
    buf g_G4679 (G4679, G1829);
    buf g_G4687 (G4687, G1704);
    buf g_G4695 (G4695, G1704);
    buf g_G4703 (G4703, G1712);
    buf g_G4711 (G4711, G1712);
    buf g_G4724 (G4724, G1749);
    not g_G4818 (G4818, G4812);
    buf g_G4855 (G4855, G1958);
    buf g_G4865 (G4865, G1966);
    buf g_G4870 (G4870, G2001);
    buf g_G4913 (G4913, G1958);
    buf g_G4923 (G4923, G1966);
    buf g_G4951 (G4951, G2106);
    buf g_G5006 (G5006, G2089);
    buf g_G5039 (G5039, G2106);
    not g_G5148 (G5148, G5142);
    not g_G5149 (G5149, G5145);
    not g_G5158 (G5158, G5152);
    not g_G5159 (G5159, G5155);
    not g_G5192 (G5192, G5186);
    not g_G5193 (G5193, G5189);
    not g_G5202 (G5202, G5196);
    not g_G5203 (G5203, G5199);
    nand g_G5284 (G5284, G5279, G5282);
    nand g_G5285 (G5285, G5276, G5283);
    nand g_G5320 (G5320, G5315, G5318);
    nand g_G5321 (G5321, G5312, G5319);
    nand g_G5386 (G5386, G5330, G5331);
    nand g_G5404 (G5404, G5399, G5402);
    and g_G598 (G598, G595, G596, G597);
    not g_G609 (G609, G3350);
    nand g_G1021 (G1021, G4119, G4122);
    nand g_G1032 (G1032, G4127, G4130);
    nand g_G1050 (G1050, G4135, G4138);
    nand g_G1078 (G1078, G4143, G4146);
    nand g_G1087 (G1087, G4151, G4154);
    nand g_G1098 (G1098, G4159, G4162);
    nand g_G1114 (G1114, G4167, G4170);
    nand g_G1132 (G1132, G4175, G4178);
    nand g_G1150 (G1150, G4183, G4186);
    nand g_G1277 (G1277, G4276, G4283);
    nand g_G1288 (G1288, G4284, G4291);
    nand g_G1306 (G1306, G4292, G4299);
    nand g_G1331 (G1331, G4300, G4307);
    nand g_G1343 (G1343, G4308, G4315);
    nand g_G1364 (G1364, G4316, G4323);
    nand g_G1389 (G1389, G4324, G4331);
    nand g_G1421 (G1421, G4332, G4339);
    nand g_G1429 (G1429, G4340, G4347);
    nand g_G1728 (G1728, G4631, G4634);
    nand g_G1756 (G1756, G4639, G4642);
    nand g_G1765 (G1765, G4647, G4650);
    nand g_G1778 (G1778, G1776, G1777);
    nand g_G1792 (G1792, G4663, G4666);
    nand g_G1810 (G1810, G4671, G4674);
    nand g_G1983 (G1983, G4764, G4771);
    nand g_G2008 (G2008, G4772, G4779);
    nand g_G2021 (G2021, G2019, G2020);
    nand g_G2041 (G2041, G4788, G4795);
    nand g_G2066 (G2066, G4796, G4803);
    nand g_G2098 (G2098, G4804, G4811);
    nand g_G3443 (G3443, G5121, G5124);
    nand g_G3444 (G3444, G5118, G5125);
    nand g_G3453 (G3453, G5126, G5133);
    nand g_G3461 (G3461, G5137, G5140);
    nand g_G3466 (G3466, G5165, G5168);
    nand g_G3467 (G3467, G5162, G5169);
    nand g_G3475 (G3475, G5173, G5176);
    nand g_G3476 (G3476, G5170, G5177);
    nand g_G3485 (G3485, G5178, G5185);
    not g_G5243 (G5243, G5239);
    nand g_G3862 (G3862, G3860, G3861);
    nand g_G3871 (G3871, G3869, G3870);
    nand g_G3883 (G3883, G3881, G3882);
    nand g_G3892 (G3892, G3890, G3891);
    nor g_G3956 (G3956, G3954, G3955);
    nor g_G3959 (G3959, G3957, G3958);
    or g_G4756 (G4756, G1837, G1875);
    nand g_G5150 (G5150, G5145, G5148);
    nand g_G5151 (G5151, G5142, G5149);
    nand g_G5160 (G5160, G5155, G5158);
    nand g_G5161 (G5161, G5152, G5159);
    nand g_G5194 (G5194, G5189, G5192);
    nand g_G5195 (G5195, G5186, G5193);
    nand g_G5204 (G5204, G5199, G5202);
    nand g_G5205 (G5205, G5196, G5203);
    nand g_G5236 (G5236, G3518, G3515);
    buf g_G5286 (G5286, G3350);
    nand g_G5379 (G5379, G5284, G5285);
    nand g_G5389 (G5389, G5320, G5321);
    nand g_G5425 (G5425, G5404, G5405);
    and g_G610 (G610, G607, G608, G609);
    nand g_G1023 (G1023, G1021, G1022);
    nand g_G1034 (G1034, G1032, G1033);
    nand g_G1052 (G1052, G1050, G1051);
    nand g_G1080 (G1080, G1078, G1079);
    nand g_G1089 (G1089, G1087, G1088);
    nand g_G1100 (G1100, G1098, G1099);
    nand g_G1116 (G1116, G1114, G1115);
    nand g_G1134 (G1134, G1132, G1133);
    nand g_G1152 (G1152, G1150, G1151);
    not g_G4242 (G4242, G4236);
    nand g_G1278 (G1278, G1276, G1277);
    nand g_G1289 (G1289, G1287, G1288);
    nand g_G1307 (G1307, G1305, G1306);
    nand g_G1332 (G1332, G1330, G1331);
    nand g_G1344 (G1344, G1342, G1343);
    nand g_G1365 (G1365, G1363, G1364);
    nand g_G1390 (G1390, G1388, G1389);
    nand g_G1422 (G1422, G1420, G1421);
    nand g_G1430 (G1430, G1428, G1429);
    nand g_G1730 (G1730, G1728, G1729);
    nand g_G1758 (G1758, G1756, G1757);
    nand g_G1767 (G1767, G1765, G1766);
    nand g_G1794 (G1794, G1792, G1793);
    nand g_G1812 (G1812, G1810, G1811);
    nand g_G1876 (G1876, G4679, G4682);
    not g_G4683 (G4683, G4679);
    not g_G4691 (G4691, G4687);
    not g_G4699 (G4699, G4695);
    not g_G4707 (G4707, G4703);
    not g_G4715 (G4715, G4711);
    not g_G4730 (G4730, G4724);
    nand g_G1984 (G1984, G1982, G1983);
    nand g_G2009 (G2009, G2007, G2008);
    nand g_G2042 (G2042, G2040, G2041);
    nand g_G2067 (G2067, G2065, G2066);
    nand g_G2099 (G2099, G2097, G2098);
    not g_G4869 (G4869, G4865);
    not g_G4927 (G4927, G4923);
    nand g_G3445 (G3445, G3443, G3444);
    nand g_G3454 (G3454, G3452, G3453);
    nand g_G3463 (G3463, G3461, G3462);
    nand g_G3468 (G3468, G3466, G3467);
    nand g_G3477 (G3477, G3475, G3476);
    nand g_G3486 (G3486, G3484, G3485);
    and g_G4103 (G4103, G4099, G3170);
    not g_G4412 (G4412, G4406);
    not g_G4558 (G4558, G4552);
    not g_G4859 (G4859, G4855);
    not g_G4876 (G4876, G4870);
    not g_G4917 (G4917, G4913);
    not g_G4955 (G4955, G4951);
    not g_G5012 (G5012, G5006);
    not g_G5043 (G5043, G5039);
    nand g_G5216 (G5216, G5160, G5161);
    nand g_G5219 (G5219, G5150, G5151);
    nand g_G5226 (G5226, G5204, G5205);
    nand g_G5229 (G5229, G5194, G5195);
    not g_G5392 (G5392, G5386);
    nand g_G5422 (G5422, G3959, G3956);
    and g_G1866 (G1866, G1778, G1806);
    nand g_G1877 (G1877, G4676, G4683);
    not g_G4762 (G4762, G4756);
    and g_G2142 (G2142, G2021, G2059);
    and g_G2146 (G2146, G2021, G2059);
    not g_G5242 (G5242, G5236);
    nand g_G3532 (G3532, G5236, G5243);
    not g_G3866 (G3866, G3862);
    not g_G3887 (G3887, G3883);
    buf g_G3918 (G3918, G3871);
    buf g_G3922 (G3922, G3871);
    buf g_G3926 (G3926, G3892);
    buf g_G3930 (G3930, G3892);
    not g_G5429 (G5429, G5425);
    or g_G4104 (G4104, G4099, G4103);
    buf g_G4743 (G4743, G1778);
    buf g_G4991 (G4991, G2021);
    buf g_G5001 (G5001, G2021);
    not g_G5292 (G5292, G5286);
    nand g_G5295 (G5295, G5286, G5293);
    not g_G5383 (G5383, G5379);
    not g_G5393 (G5393, G5389);
    nand g_G5394 (G5394, G5389, G5392);
    and g_G1439 (G1439, G1278, G1301);
    and g_G1440 (G1440, G1289, G1278, G1318);
    and g_G1441 (G1441, G1307, G1278, G1324, G1289);
    and g_G1847 (G1847, G1730, G1704, G1749, G1712);
    and g_G1168 (G1168, G1023, G1046);
    and g_G1169 (G1169, G1034, G1023, G1064);
    and g_G1170 (G1170, G1052, G1023, G1071, G1034);
    and g_G2117 (G2117, G1984, G1958, G2001, G1966);
    not g_G1086 (G1086, G1080);
    and g_G1166 (G1166, G1034, G1080, G1052, G1023);
    and g_G1171 (G1171, G1034, G1064);
    and g_G1172 (G1172, G1052, G1071, G1034);
    and g_G1173 (G1173, G1080, G1052, G1034);
    and g_G1174 (G1174, G1034, G1064);
    and g_G1175 (G1175, G1071, G1052, G1034);
    and g_G1176 (G1176, G1052, G1071);
    and g_G1177 (G1177, G1080, G1052);
    and g_G1178 (G1178, G1052, G1071);
    and g_G1179 (G1179, G1100, G1179_tmp);
    and g_G1179_tmp (G1179_tmp, G1152, G1116, G1089, G1134);
    and g_G1181 (G1181, G1089, G1111);
    and g_G1182 (G1182, G1100, G1089, G1128);
    and g_G1183 (G1183, G1116, G1089, G1145, G1100);
    and g_G1184 (G1184, G1134, G1184_tmp);
    and g_G1184_tmp (G1184_tmp, G1116, G1089, G1160, G1100);
    and g_G1188 (G1188, G1100, G1128);
    and g_G1189 (G1189, G1116, G1145, G1100);
    and g_G1190 (G1190, G1134, G1116, G1160, G1100);
    and g_G1191 (G1191, G4, G1191_tmp);
    and g_G1191_tmp (G1191_tmp, G1152, G1116, G1134, G1100);
    and g_G1192 (G1192, G1145, G1116);
    and g_G1193 (G1193, G1134, G1116, G1160);
    and g_G1194 (G1194, G4, G1152, G1116, G1134);
    and g_G1195 (G1195, G1134, G1160);
    and g_G1196 (G1196, G4, G1152, G1134);
    and g_G1197 (G1197, G4, G1152);
    and g_G1437 (G1437, G1422, G1307, G1289, G1278);
    and g_G1442 (G1442, G1289, G1318);
    and g_G1443 (G1443, G1307, G1324, G1289);
    and g_G1444 (G1444, G1422, G1307, G1289);
    and g_G1445 (G1445, G1289, G1318);
    and g_G1446 (G1446, G1307, G1324, G1289);
    and g_G1447 (G1447, G1307, G1324);
    and g_G1451 (G1451, G1430, G1451_tmp);
    and g_G1451_tmp (G1451_tmp, G1390, G1365, G1344, G1332);
    and g_G1454 (G1454, G1332, G1359);
    and g_G1455 (G1455, G1344, G1332, G1382);
    and g_G1456 (G1456, G1365, G1332, G1404, G1344);
    and g_G1457 (G1457, G1390, G1457_tmp);
    and g_G1457_tmp (G1457_tmp, G1365, G1332, G1412, G1344);
    and g_G1465 (G1465, G1344, G1382);
    and g_G1466 (G1466, G1365, G1404, G1344);
    and g_G1467 (G1467, G1390, G1365, G1412, G1344);
    and g_G1468 (G1468, G1430, G1365, G1344, G1390);
    and g_G1469 (G1469, G1344, G1382);
    and g_G1470 (G1470, G1365, G1404, G1344);
    and g_G1471 (G1471, G1390, G1365, G1412, G1344);
    and g_G1472 (G1472, G1365, G1404);
    and g_G1473 (G1473, G1390, G1365, G1412);
    and g_G1474 (G1474, G1430, G1365, G1390);
    and g_G1475 (G1475, G1365, G1404);
    and g_G1476 (G1476, G1390, G1365, G1412);
    and g_G1477 (G1477, G1390, G1412);
    and g_G1481 (G1481, G1422, G1307);
    and g_G1482 (G1482, G1430, G1390);
    not g_G1764 (G1764, G1758);
    and g_G1843 (G1843, G1712, G1758, G1730, G1704);
    and g_G1850 (G1850, G1730, G1749, G1712);
    and g_G1851 (G1851, G1758, G1730, G1712);
    and g_G1853 (G1853, G1749, G1730, G1712);
    and g_G1854 (G1854, G1730, G1749);
    and g_G1855 (G1855, G1758, G1730);
    and g_G1856 (G1856, G1730, G1749);
    and g_G1857 (G1857, G1778, G1857_tmp);
    and g_G1857_tmp (G1857_tmp, G1829, G1794, G1767, G1812);
    and g_G1859 (G1859, G1767, G1789);
    and g_G1860 (G1860, G1778, G1767, G1806);
    and g_G1861 (G1861, G1794, G1767, G1823, G1778);
    and g_G1862 (G1862, G1812, G1862_tmp);
    and g_G1862_tmp (G1862_tmp, G1794, G1767, G1837, G1778);
    and g_G1867 (G1867, G1794, G1823, G1778);
    and g_G1868 (G1868, G1812, G1794, G1837, G1778);
    and g_G1869 (G1869, G54, G1869_tmp);
    and g_G1869_tmp (G1869_tmp, G1829, G1794, G1812, G1778);
    and g_G1870 (G1870, G1823, G1794);
    and g_G1871 (G1871, G1812, G1794, G1837);
    and g_G1872 (G1872, G54, G1829, G1794, G1812);
    and g_G1873 (G1873, G1812, G1837);
    and g_G1874 (G1874, G54, G1829, G1812);
    nand g_G1878 (G1878, G1876, G1877);
    and g_G2113 (G2113, G2099, G1984, G1966, G1958);
    and g_G2120 (G2120, G1984, G2001, G1966);
    and g_G2121 (G2121, G2099, G1984, G1966);
    and g_G2123 (G2123, G1984, G2001, G1966);
    and g_G2124 (G2124, G1984, G2001);
    and g_G2128 (G2128, G2106, G2128_tmp);
    and g_G2128_tmp (G2128_tmp, G2067, G2042, G2021, G2009);
    and g_G2131 (G2131, G2009, G2036);
    and g_G2132 (G2132, G2021, G2009, G2059);
    and g_G2133 (G2133, G2042, G2009, G2081, G2021);
    and g_G2134 (G2134, G2067, G2134_tmp);
    and g_G2134_tmp (G2134_tmp, G2042, G2009, G2089, G2021);
    and g_G2143 (G2143, G2042, G2081, G2021);
    and g_G2144 (G2144, G2067, G2042, G2089, G2021);
    and g_G2145 (G2145, G2106, G2042, G2021, G2067);
    and g_G2147 (G2147, G2042, G2081, G2021);
    and g_G2148 (G2148, G2067, G2042, G2089, G2021);
    and g_G2149 (G2149, G2042, G2081);
    and g_G2150 (G2150, G2067, G2042, G2089);
    and g_G2151 (G2151, G2106, G2042, G2067);
    and g_G2152 (G2152, G2042, G2081);
    and g_G2153 (G2153, G2067, G2042, G2089);
    and g_G2154 (G2154, G2067, G2089);
    and g_G2158 (G2158, G2099, G1984);
    and g_G2159 (G2159, G2106, G2067);
    not g_G3449 (G3449, G3445);
    not g_G3458 (G3458, G3454);
    not g_G3472 (G3472, G3468);
    not g_G3481 (G3481, G3477);
    buf g_G3497 (G3497, G3463);
    buf g_G3501 (G3501, G3463);
    buf g_G3505 (G3505, G3486);
    buf g_G3509 (G3509, G3486);
    nand g_G3531 (G3531, G5239, G5242);
    not g_G5428 (G5428, G5422);
    nand g_G3967 (G3967, G5422, G5429);
    buf g_G4191 (G4191, G1152);
    buf g_G4199 (G4199, G1023);
    buf g_G4207 (G4207, G1023);
    buf g_G4215 (G4215, G1034);
    buf g_G4223 (G4223, G1034);
    buf g_G4231 (G4231, G1052);
    buf g_G4239 (G4239, G1052);
    buf g_G4247 (G4247, G1089);
    buf g_G4255 (G4255, G1100);
    buf g_G4263 (G4263, G1116);
    buf g_G4271 (G4271, G1134);
    buf g_G4371 (G4371, G1422);
    buf g_G4381 (G4381, G1307);
    buf g_G4391 (G4391, G1278);
    buf g_G4401 (G4401, G1289);
    buf g_G4429 (G4429, G1422);
    buf g_G4439 (G4439, G1307);
    buf g_G4449 (G4449, G1278);
    buf g_G4459 (G4459, G1289);
    buf g_G4497 (G4497, G1430);
    buf g_G4507 (G4507, G1390);
    buf g_G4517 (G4517, G1332);
    buf g_G4527 (G4527, G1365);
    buf g_G4537 (G4537, G1344);
    buf g_G4547 (G4547, G1344);
    buf g_G4585 (G4585, G1430);
    buf g_G4595 (G4595, G1390);
    buf g_G4605 (G4605, G1332);
    buf g_G4615 (G4615, G1365);
    buf g_G4719 (G4719, G1730);
    buf g_G4727 (G4727, G1730);
    buf g_G4735 (G4735, G1767);
    buf g_G4751 (G4751, G1794);
    buf g_G4759 (G4759, G1812);
    buf g_G4835 (G4835, G2099);
    buf g_G4845 (G4845, G1984);
    buf g_G4893 (G4893, G2099);
    buf g_G4903 (G4903, G1984);
    buf g_G4961 (G4961, G2067);
    buf g_G4971 (G4971, G2009);
    buf g_G4981 (G4981, G2042);
    buf g_G5049 (G5049, G2067);
    buf g_G5059 (G5059, G2009);
    buf g_G5069 (G5069, G2042);
    not g_G5222 (G5222, G5216);
    not g_G5223 (G5223, G5219);
    not g_G5232 (G5232, G5226);
    not g_G5233 (G5233, G5229);
    nand g_G5294 (G5294, G5289, G5292);
    nand g_G5395 (G5395, G5386, G5393);
    or g_G589 (G589, G1286, G1439, G1440, G1441);
    or g_G616 (G616, G3167, G1845, G1846, G1847);
    or g_G619 (G619, G1031, G1168, G1169, G1170);
    or g_G627 (G627, G3167, G2115, G2116, G2117);
    or g_G1185 (G1185, G1097, G1185_tmp);
    or g_G1185_tmp (G1185_tmp, G1181, G1182, G1183, G1184);
    or g_G1448 (G1448, G1318, G1447);
    or g_G1458 (G1458, G1341, G1458_tmp);
    or g_G1458_tmp (G1458_tmp, G1454, G1455, G1456, G1457);
    or g_G1478 (G1478, G1404, G1477);
    or g_G1863 (G1863, G1775, G1863_tmp);
    or g_G1863_tmp (G1863_tmp, G1859, G1860, G1861, G1862);
    not g_G4747 (G4747, G4743);
    or g_G2125 (G2125, G1995, G2124);
    or g_G2135 (G2135, G2018, G2135_tmp);
    or g_G2135_tmp (G2135_tmp, G2131, G2132, G2133, G2134);
    or g_G2155 (G2155, G2081, G2154);
    not g_G4995 (G4995, G4991);
    not g_G5005 (G5005, G5001);
    nand g_G3533 (G3533, G3531, G3532);
    not g_G3921 (G3921, G3918);
    not g_G3925 (G3925, G3922);
    not g_G3929 (G3929, G3926);
    not g_G3933 (G3933, G3930);
    and g_G3943 (G3943, G3862, G3853, G3918);
    and g_G3946 (G3946, G3866, G3857, G3922);
    and g_G3949 (G3949, G3883, G3874, G3926);
    and g_G3952 (G3952, G3887, G3878, G3930);
    nand g_G3966 (G3966, G5425, G5428);
    nand g_G4107 (G4107, G4104, G132);
    or g_G4196 (G4196, G1046, G1171, G1172, G1173);
    nor g_G4204 (G4204, G1046, G1174, G1175);
    or g_G4212 (G4212, G1064, G1176, G1177);
    nor g_G4220 (G4220, G1064, G1178);
    or g_G4244 (G4244, G1111, G4244_tmp);
    or g_G4244_tmp (G4244_tmp, G1188, G1189, G1190, G1191);
    or g_G4252 (G4252, G1128, G1192, G1193, G1194);
    or g_G4260 (G4260, G1145, G1195, G1196);
    or g_G4268 (G4268, G1160, G1197);
    or g_G4361 (G4361, G1301, G1442, G1443, G1444);
    nor g_G4419 (G4419, G1301, G1445, G1446);
    or g_G4467 (G4467, G1382, G1472, G1473, G1474);
    or g_G4487 (G4487, G1359, G4487_tmp);
    or g_G4487_tmp (G4487_tmp, G1465, G1466, G1467, G1468);
    nor g_G4555 (G4555, G1382, G1475, G1476);
    nor g_G4575 (G4575, G1359, G1469, G1470, G1471);
    or g_G4684 (G4684, G1724, G1849, G1850, G1851);
    nor g_G4692 (G4692, G1724, G1852, G1853);
    or g_G4700 (G4700, G1742, G1854, G1855);
    nor g_G4708 (G4708, G1742, G1856);
    or g_G4732 (G4732, G1789, G4732_tmp);
    or g_G4732_tmp (G4732_tmp, G1866, G1867, G1868, G1869);
    or g_G4740 (G4740, G1806, G1870, G1871, G1872);
    or g_G4748 (G4748, G1823, G1873, G1874);
    or g_G4825 (G4825, G1978, G2119, G2120, G2121);
    nor g_G4883 (G4883, G1978, G2122, G2123);
    or g_G4928 (G4928, G2059, G2149, G2150, G2151);
    or g_G4941 (G4941, G2036, G4941_tmp);
    or g_G4941_tmp (G4941_tmp, G2142, G2143, G2144, G2145);
    nor g_G5009 (G5009, G2059, G2152, G2153);
    nor g_G5029 (G5029, G2036, G2146, G2147, G2148);
    nand g_G5224 (G5224, G5219, G5222);
    nand g_G5225 (G5225, G5216, G5223);
    nand g_G5234 (G5234, G5229, G5232);
    nand g_G5235 (G5235, G5226, G5233);
    nand g_G5376 (G5376, G5294, G5295);
    nand g_G5417 (G5417, G5394, G5395);
    not g_G576 (G576, G1878);
    and g_G588 (G588, G1437, G1451);
    and g_G615 (G615, G1843, G1857);
    and g_G626 (G626, G2113, G2128);
    and g_G632 (G632, G1166, G1179);
    nand g_G1198 (G1198, G4191, G4194);
    not g_G4195 (G4195, G4191);
    not g_G4203 (G4203, G4199);
    not g_G4211 (G4211, G4207);
    not g_G4219 (G4219, G4215);
    not g_G4227 (G4227, G4223);
    nand g_G1217 (G1217, G4231, G4234);
    not g_G4235 (G4235, G4231);
    nand g_G1221 (G1221, G4239, G4242);
    not g_G4243 (G4243, G4239);
    and g_G1224 (G1224, G1179, G4);
    not g_G4251 (G4251, G4247);
    not g_G4259 (G4259, G4255);
    not g_G4267 (G4267, G4263);
    not g_G4275 (G4275, G4271);
    not g_G1453 (G1453, G1451);
    not g_G4405 (G4405, G4401);
    not g_G4463 (G4463, G4459);
    not g_G4541 (G4541, G4537);
    not g_G4551 (G4551, G4547);
    nand g_G1895 (G1895, G4719, G4722);
    not g_G4723 (G4723, G4719);
    nand g_G1899 (G1899, G4727, G4730);
    not g_G4731 (G4731, G4727);
    and g_G1902 (G1902, G1857, G54);
    not g_G4739 (G4739, G4735);
    not g_G4755 (G4755, G4751);
    nand g_G1929 (G1929, G4759, G4762);
    not g_G4763 (G4763, G4759);
    not g_G2130 (G2130, G2128);
    not g_G3500 (G3500, G3497);
    not g_G3504 (G3504, G3501);
    not g_G3508 (G3508, G3505);
    not g_G3512 (G3512, G3509);
    and g_G3520 (G3520, G3454, G3445, G3497);
    and g_G3523 (G3523, G3458, G3449, G3501);
    and g_G3526 (G3526, G3477, G3468, G3505);
    and g_G3529 (G3529, G3481, G3472, G3509);
    buf g_G1002 (G1002, G3533);
    and g_G3837 (G3837, G1878, G3795, G3823);
    and g_G3942 (G3942, G3857, G3862, G3921);
    and g_G3945 (G3945, G3853, G3866, G3925);
    and g_G3948 (G3948, G3878, G3883, G3929);
    and g_G3951 (G3951, G3874, G3887, G3933);
    nand g_G3968 (G3968, G3966, G3967);
    not g_G4375 (G4375, G4371);
    not g_G4385 (G4385, G4381);
    not g_G4395 (G4395, G4391);
    not g_G4433 (G4433, G4429);
    not g_G4443 (G4443, G4439);
    not g_G4453 (G4453, G4449);
    not g_G4501 (G4501, G4497);
    not g_G4511 (G4511, G4507);
    not g_G4521 (G4521, G4517);
    not g_G4531 (G4531, G4527);
    not g_G4619 (G4619, G4615);
    not g_G4589 (G4589, G4585);
    not g_G4599 (G4599, G4595);
    not g_G4609 (G4609, G4605);
    not g_G4839 (G4839, G4835);
    not g_G4849 (G4849, G4845);
    not g_G4897 (G4897, G4893);
    not g_G4907 (G4907, G4903);
    not g_G4965 (G4965, G4961);
    not g_G4975 (G4975, G4971);
    not g_G4985 (G4985, G4981);
    not g_G5073 (G5073, G5069);
    not g_G5053 (G5053, G5049);
    not g_G5063 (G5063, G5059);
    nand g_G5247 (G5247, G5224, G5225);
    nand g_G5255 (G5255, G5234, G5235);
    and g_G590 (G590, G1437, G1458);
    and g_G617 (G617, G1863, G1843);
    and g_G620 (G620, G1185, G1166);
    and g_G628 (G628, G2113, G2135);
    not g_G3535 (G3535, G3533);
    nand g_G1199 (G1199, G4188, G4195);
    not g_G4202 (G4202, G4196);
    nand g_G1204 (G1204, G4196, G4203);
    not g_G4210 (G4210, G4204);
    nand g_G1207 (G1207, G4204, G4211);
    not g_G4218 (G4218, G4212);
    nand g_G1211 (G1211, G4212, G4219);
    not g_G4226 (G4226, G4220);
    nand g_G1214 (G1214, G4220, G4227);
    nand g_G1218 (G1218, G4228, G4235);
    nand g_G1222 (G1222, G4236, G4243);
    or g_G1225 (G1225, G1185, G1224);
    not g_G4250 (G4250, G4244);
    nand g_G1237 (G1237, G4244, G4251);
    not g_G4258 (G4258, G4252);
    nand g_G1242 (G1242, G4252, G4259);
    not g_G4266 (G4266, G4260);
    nand g_G1247 (G1247, G4260, G4267);
    not g_G4274 (G4274, G4268);
    nand g_G1252 (G1252, G4268, G4275);
    not g_G1462 (G1462, G1458);
    not g_G4690 (G4690, G4684);
    nand g_G1882 (G1882, G4684, G4691);
    not g_G4698 (G4698, G4692);
    nand g_G1885 (G1885, G4692, G4699);
    not g_G4706 (G4706, G4700);
    nand g_G1889 (G1889, G4700, G4707);
    not g_G4714 (G4714, G4708);
    nand g_G1892 (G1892, G4708, G4715);
    nand g_G1896 (G1896, G4716, G4723);
    nand g_G1900 (G1900, G4724, G4731);
    or g_G1903 (G1903, G1863, G1902);
    not g_G4738 (G4738, G4732);
    nand g_G1915 (G1915, G4732, G4739);
    not g_G4746 (G4746, G4740);
    nand g_G1920 (G1920, G4740, G4747);
    not g_G4754 (G4754, G4748);
    nand g_G1925 (G1925, G4748, G4755);
    nand g_G1930 (G1930, G4756, G4763);
    not g_G2139 (G2139, G2135);
    and g_G3519 (G3519, G3449, G3454, G3500);
    and g_G3522 (G3522, G3445, G3458, G3504);
    and g_G3525 (G3525, G3472, G3477, G3508);
    and g_G3528 (G3528, G3468, G3481, G3512);
    or g_G3848 (G3848, G3836, G3837, G3838);
    nor g_G3944 (G3944, G3942, G3943);
    nor g_G3947 (G3947, G3945, G3946);
    nor g_G3950 (G3950, G3948, G3949);
    nor g_G3953 (G3953, G3951, G3952);
    not g_G5421 (G5421, G5417);
    buf g_G1004 (G1004, G3968);
    and g_G4111 (G4111, G4104, G4107);
    and g_G4112 (G4112, G4107, G132);
    or g_G4351 (G4351, G1448, G1481);
    not g_G4365 (G4365, G4361);
    not g_G4409 (G4409, G1448);
    not g_G4423 (G4423, G4419);
    not g_G4471 (G4471, G4467);
    nand g_G4472 (G4472, G4467, G4470);
    or g_G4477 (G4477, G1478, G1482);
    not g_G4491 (G4491, G4487);
    not g_G4559 (G4559, G4555);
    nand g_G4560 (G4560, G4555, G4558);
    not g_G4565 (G4565, G1478);
    not g_G4579 (G4579, G4575);
    or g_G4815 (G4815, G2125, G2158);
    not g_G4829 (G4829, G4825);
    not g_G4873 (G4873, G2125);
    not g_G4887 (G4887, G4883);
    or g_G4931 (G4931, G2155, G2159);
    not g_G4934 (G4934, G4928);
    not g_G4945 (G4945, G4941);
    not g_G5013 (G5013, G5009);
    nand g_G5014 (G5014, G5009, G5012);
    not g_G5019 (G5019, G2155);
    not g_G5033 (G5033, G5029);
    not g_G5382 (G5382, G5376);
    nand g_G5385 (G5385, G5376, G5383);
    or g_G591 (G591, G589, G590);
    or g_G618 (G618, G616, G617);
    or g_G621 (G621, G619, G620);
    or g_G629 (G629, G627, G628);
    not g_G3970 (G3970, G3968);
    nand g_G1200 (G1200, G1198, G1199);
    nand g_G1203 (G1203, G4199, G4202);
    nand g_G1206 (G1206, G4207, G4210);
    nand g_G1210 (G1210, G4215, G4218);
    nand g_G1213 (G1213, G4223, G4226);
    nand g_G1219 (G1219, G1217, G1218);
    nand g_G1223 (G1223, G1221, G1222);
    nand g_G1236 (G1236, G4247, G4250);
    nand g_G1241 (G1241, G4255, G4258);
    nand g_G1246 (G1246, G4263, G4266);
    nand g_G1251 (G1251, G4271, G4274);
    nand g_G1881 (G1881, G4687, G4690);
    nand g_G1884 (G1884, G4695, G4698);
    nand g_G1888 (G1888, G4703, G4706);
    nand g_G1891 (G1891, G4711, G4714);
    nand g_G1897 (G1897, G1895, G1896);
    nand g_G1901 (G1901, G1899, G1900);
    nand g_G1914 (G1914, G4735, G4738);
    nand g_G1919 (G1919, G4743, G4746);
    nand g_G1924 (G1924, G4751, G4754);
    nand g_G1931 (G1931, G1929, G1930);
    nor g_G3521 (G3521, G3519, G3520);
    nor g_G3524 (G3524, G3522, G3523);
    nor g_G3527 (G3527, G3525, G3526);
    nor g_G3530 (G3530, G3528, G3529);
    not g_G5251 (G5251, G5247);
    not g_G5259 (G5259, G5255);
    or g_G4113 (G4113, G4111, G4112);
    nand g_G4473 (G4473, G4464, G4471);
    nand g_G4561 (G4561, G4552, G4559);
    nand g_G5015 (G5015, G5006, G5013);
    nand g_G5384 (G5384, G5379, G5382);
    nand g_G5406 (G5406, G3947, G3944);
    nand g_G5414 (G5414, G3953, G3950);
    and g_G1664 (G1664, G3848, G1621, G1645);
    and g_G2335 (G2335, G3848, G2293, G2316);
    and g_G718 (G718, G3848, G2430, G2454);
    not g_G822 (G822, G3848);
    and g_G855 (G855, G3848, G2488, G2512);
    nand g_G1205 (G1205, G1203, G1204);
    nand g_G1208 (G1208, G1206, G1207);
    nand g_G1212 (G1212, G1210, G1211);
    nand g_G1215 (G1215, G1213, G1214);
    not g_G1220 (G1220, G1219);
    not g_G1231 (G1231, G1225);
    nand g_G1238 (G1238, G1236, G1237);
    nand g_G1243 (G1243, G1241, G1242);
    nand g_G1248 (G1248, G1246, G1247);
    nand g_G1253 (G1253, G1251, G1252);
    and g_G1272 (G1272, G1225, G1086);
    and g_G1483 (G1483, G1462, G1453);
    nand g_G1883 (G1883, G1881, G1882);
    nand g_G1886 (G1886, G1884, G1885);
    nand g_G1890 (G1890, G1888, G1889);
    nand g_G1893 (G1893, G1891, G1892);
    not g_G1898 (G1898, G1897);
    not g_G1909 (G1909, G1903);
    nand g_G1916 (G1916, G1914, G1915);
    nand g_G1921 (G1921, G1919, G1920);
    nand g_G1926 (G1926, G1924, G1925);
    and g_G1953 (G1953, G1903, G1764);
    and g_G2160 (G2160, G2139, G2130);
    not g_G4355 (G4355, G4351);
    nand g_G4356 (G4356, G4351, G4354);
    not g_G4413 (G4413, G4409);
    nand g_G4414 (G4414, G4409, G4412);
    nand g_G4474 (G4474, G4472, G4473);
    not g_G4481 (G4481, G4477);
    nand g_G4562 (G4562, G4560, G4561);
    not g_G4569 (G4569, G4565);
    not g_G4819 (G4819, G4815);
    nand g_G4820 (G4820, G4815, G4818);
    not g_G4877 (G4877, G4873);
    nand g_G4878 (G4878, G4873, G4876);
    not g_G4935 (G4935, G4931);
    nand g_G4936 (G4936, G4931, G4934);
    nand g_G5016 (G5016, G5014, G5015);
    not g_G5023 (G5023, G5019);
    nand g_G5244 (G5244, G3524, G3521);
    nand g_G5252 (G5252, G3530, G3527);
    nand g_G5409 (G5409, G5384, G5385);
    not g_G566 (G566, G1200);
    not g_G577 (G577, G1931);
    and g_G3733 (G3733, G4113, G3724, G3721);
    not g_G1209 (G1209, G1208);
    not g_G1216 (G1216, G1215);
    and g_G1257 (G1257, G1225, G1205);
    and g_G1262 (G1262, G1225, G1212);
    and g_G1267 (G1267, G1225, G1220);
    not g_G1887 (G1887, G1886);
    not g_G1894 (G1894, G1893);
    and g_G1935 (G1935, G1903, G1883);
    and g_G1943 (G1943, G1903, G1890);
    and g_G1948 (G1948, G1903, G1898);
    and g_G3779 (G3779, G1200, G3737, G3765);
    and g_G3840 (G3840, G1931, G3795, G3823);
    not g_G5412 (G5412, G5406);
    not g_G5420 (G5420, G5414);
    nand g_G3964 (G3964, G5414, G5421);
    nand g_G4357 (G4357, G4348, G4355);
    nand g_G4415 (G4415, G4406, G4413);
    nand g_G4821 (G4821, G4812, G4819);
    nand g_G4879 (G4879, G4870, G4877);
    nand g_G4937 (G4937, G4928, G4935);
    not g_G567 (G567, G1253);
    not g_G568 (G568, G1248);
    not g_G569 (G569, G1243);
    not g_G570 (G570, G1238);
    not g_G578 (G578, G1926);
    not g_G579 (G579, G1921);
    not g_G580 (G580, G1916);
    and g_G1256 (G1256, G1209, G1231);
    and g_G1261 (G1261, G1216, G1231);
    and g_G1266 (G1266, G1223, G1231);
    and g_G1271 (G1271, G1080, G1231);
    not g_G1486 (G1486, G1483);
    and g_G1934 (G1934, G1887, G1909);
    and g_G1942 (G1942, G1894, G1909);
    and g_G1947 (G1947, G1901, G1909);
    and g_G1952 (G1952, G1758, G1909);
    not g_G2163 (G2163, G2160);
    not g_G5250 (G5250, G5244);
    nand g_G3537 (G3537, G5244, G5251);
    not g_G5258 (G5258, G5252);
    nand g_G3542 (G3542, G5252, G5259);
    and g_G3782 (G3782, G1253, G3737, G3765);
    and g_G3785 (G3785, G1248, G3737, G3765);
    and g_G3788 (G3788, G1243, G3737, G3765);
    or g_G3790 (G3790, G3778, G3779, G3780);
    and g_G3843 (G3843, G1926, G3795, G3823);
    and g_G3846 (G3846, G1921, G3795, G3823);
    or g_G3849 (G3849, G3839, G3840, G3841);
    nand g_G3960 (G3960, G5409, G5412);
    not g_G5413 (G5413, G5409);
    nand g_G3963 (G3963, G5417, G5420);
    and g_G4010 (G4010, G1238, G3972, G3998);
    and g_G4068 (G4068, G1916, G4030, G4056);
    nand g_G4358 (G4358, G4356, G4357);
    nand g_G4416 (G4416, G4414, G4415);
    not g_G4480 (G4480, G4474);
    nand g_G4483 (G4483, G4474, G4481);
    not g_G4568 (G4568, G4562);
    nand g_G4571 (G4571, G4562, G4569);
    nand g_G4822 (G4822, G4820, G4821);
    nand g_G4880 (G4880, G4878, G4879);
    nand g_G4938 (G4938, G4936, G4937);
    not g_G5022 (G5022, G5016);
    nand g_G5025 (G5025, G5016, G5023);
    or g_G1258 (G1258, G1256, G1257);
    or g_G1263 (G1263, G1261, G1262);
    or g_G1268 (G1268, G1266, G1267);
    or g_G1273 (G1273, G1271, G1272);
    or g_G1936 (G1936, G1934, G1935);
    or g_G1944 (G1944, G1942, G1943);
    or g_G1949 (G1949, G1947, G1948);
    or g_G1954 (G1954, G1952, G1953);
    nand g_G3536 (G3536, G5247, G5250);
    nand g_G3541 (G3541, G5255, G5258);
    or g_G3791 (G3791, G3781, G3782, G3783);
    or g_G3792 (G3792, G3784, G3785, G3786);
    or g_G3793 (G3793, G3787, G3788, G3789);
    or g_G3850 (G3850, G3842, G3843, G3844);
    or g_G3851 (G3851, G3845, G3846, G3847);
    nand g_G3961 (G3961, G5406, G5413);
    nand g_G3965 (G3965, G3963, G3964);
    or g_G4024 (G4024, G4009, G4010, G4011);
    or g_G4082 (G4082, G4067, G4068, G4069);
    nand g_G4482 (G4482, G4477, G4480);
    nand g_G4570 (G4570, G4565, G4568);
    nand g_G5024 (G5024, G5019, G5022);
    and g_G1666 (G1666, G3790, G1609, G1645);
    and g_G1670 (G1670, G3849, G1621, G1645);
    and g_G2337 (G2337, G3790, G2281, G2316);
    and g_G2341 (G2341, G3849, G2293, G2316);
    and g_G719 (G719, G3790, G2418, G2454);
    and g_G758 (G758, G3849, G2430, G2454);
    and g_G798 (G798, G3849, G2488, G2512);
    not g_G838 (G838, G3849);
    and g_G856 (G856, G3790, G2476, G2512);
    not g_G861 (G861, G3790);
    nand g_G3538 (G3538, G3536, G3537);
    nand g_G3543 (G3543, G3541, G3542);
    nand g_G3962 (G3962, G3960, G3961);
    not g_G4364 (G4364, G4358);
    nand g_G4367 (G4367, G4358, G4365);
    not g_G4422 (G4422, G4416);
    nand g_G4425 (G4425, G4416, G4423);
    nand g_G4484 (G4484, G4482, G4483);
    nand g_G4572 (G4572, G4570, G4571);
    not g_G4828 (G4828, G4822);
    nand g_G4831 (G4831, G4822, G4829);
    not g_G4886 (G4886, G4880);
    nand g_G4889 (G4889, G4880, G4887);
    not g_G4944 (G4944, G4938);
    nand g_G4947 (G4947, G4938, G4945);
    nand g_G5026 (G5026, G5024, G5025);
    not g_G571 (G571, G1273);
    not g_G572 (G572, G1268);
    not g_G573 (G573, G1263);
    not g_G574 (G574, G1258);
    not g_G581 (G581, G1954);
    not g_G582 (G582, G1949);
    not g_G583 (G583, G1944);
    not g_G584 (G584, G1936);
    not g_G623 (G623, G1936);
    and g_G1576 (G1576, G4082, G1540, G1564);
    and g_G1578 (G1578, G4024, G1528, G1564);
    or g_G659 (G659, G1664, G1666, G1667, G1668);
    and g_G1672 (G1672, G3791, G1609, G1645);
    and g_G1676 (G1676, G3850, G1621, G1645);
    and g_G1678 (G1678, G3792, G1609, G1645);
    and g_G1682 (G1682, G3851, G1621, G1645);
    and g_G1684 (G1684, G3793, G1609, G1645);
    and g_G2250 (G2250, G4082, G2215, G2238);
    and g_G2252 (G2252, G4024, G2203, G2238);
    or g_G691 (G691, G2335, G2337, G2338, G2339);
    and g_G2343 (G2343, G3791, G2281, G2316);
    and g_G2347 (G2347, G3850, G2293, G2316);
    and g_G2349 (G2349, G3792, G2281, G2316);
    and g_G2353 (G2353, G3851, G2293, G2316);
    and g_G2355 (G2355, G3793, G2281, G2316);
    or g_G722 (G722, G718, G719, G720, G721);
    and g_G743 (G743, G4082, G3570, G3594);
    and g_G744 (G744, G4024, G3558, G3594);
    and g_G748 (G748, G3851, G2430, G2454);
    and g_G749 (G749, G3793, G2418, G2454);
    and g_G753 (G753, G3850, G2430, G2454);
    and g_G754 (G754, G3792, G2418, G2454);
    and g_G759 (G759, G3791, G2418, G2454);
    and g_G783 (G783, G4082, G3672, G3696);
    and g_G784 (G784, G4024, G3660, G3696);
    and g_G788 (G788, G3851, G2488, G2512);
    and g_G789 (G789, G3793, G2476, G2512);
    and g_G793 (G793, G3850, G2488, G2512);
    and g_G794 (G794, G3792, G2476, G2512);
    and g_G799 (G799, G3791, G2476, G2512);
    and g_G3735 (G3735, G1936, G3724, G3717);
    not g_G832 (G832, G4082);
    not g_G834 (G834, G3851);
    not g_G836 (G836, G3850);
    not g_G3835 (G3835, G3965);
    or g_G859 (G859, G855, G856, G857, G858);
    not g_G871 (G871, G4024);
    not g_G873 (G873, G3793);
    not g_G875 (G875, G3792);
    not g_G877 (G877, G3791);
    buf g_G998 (G998, G3538);
    buf g_G1000 (G1000, G3543);
    and g_G3651 (G3651, G3965, G3632);
    and g_G4013 (G4013, G1273, G3972, G3998);
    and g_G4016 (G4016, G1268, G3972, G3998);
    and g_G4019 (G4019, G1263, G3972, G3998);
    and g_G4022 (G4022, G1258, G3972, G3998);
    and g_G4071 (G4071, G1954, G4030, G4056);
    and g_G4074 (G4074, G1949, G4030, G4056);
    and g_G4077 (G4077, G1944, G4030, G4056);
    and g_G4080 (G4080, G1936, G4030, G4056);
    nand g_G4096 (G4096, G4113, G1936);
    nand g_G4366 (G4366, G4361, G4364);
    nand g_G4424 (G4424, G4419, G4422);
    nand g_G4830 (G4830, G4825, G4828);
    nand g_G4888 (G4888, G4883, G4886);
    nand g_G4946 (G4946, G4941, G4944);
    and g_G575 (G575, G566, G575_0_tmp, G575_1_tmp);
    and g_G575_0_tmp (G575_0_tmp, G567, G568, G569, G570);
    and g_G575_1_tmp (G575_1_tmp, G571, G572, G573, G574);
    and g_G585 (G585, G576, G585_0_tmp, G585_1_tmp);
    and g_G585_0_tmp (G585_0_tmp, G577, G578, G579, G580);
    and g_G585_1_tmp (G585_1_tmp, G581, G582, G583, G584);
    or g_G640 (G640, G1576, G1578, G1579, G1580);
    and g_G661 (G661, G659, G1606);
    or g_G662 (G662, G1670, G1672, G1673, G1674);
    or g_G665 (G665, G1676, G1678, G1679, G1680);
    or g_G668 (G668, G1682, G1684, G1685, G1686);
    or g_G674 (G674, G2250, G2252, G2253, G2254);
    and g_G693 (G693, G691, G2279);
    or g_G694 (G694, G2341, G2343, G2344, G2345);
    or g_G697 (G697, G2347, G2349, G2350, G2351);
    or g_G700 (G700, G2353, G2355, G2356, G2357);
    or g_G747 (G747, G743, G744, G745, G746);
    or g_G752 (G752, G748, G749, G750, G751);
    or g_G757 (G757, G753, G754, G755, G756);
    or g_G762 (G762, G758, G759, G760, G761);
    or g_G787 (G787, G783, G784, G785, G786);
    or g_G792 (G792, G788, G789, G790, G791);
    or g_G797 (G797, G793, G794, G795, G796);
    or g_G802 (G802, G798, G799, G800, G801);
    or g_G817 (G817, G3731, G3733, G3734, G3735);
    and g_G839 (G839, G3835, G3803, G3823);
    not g_G3540 (G3540, G3538);
    not g_G3545 (G3545, G3543);
    not g_G3777 (G3777, G3962);
    and g_G3648 (G3648, G3962, G3632);
    or g_G4025 (G4025, G4012, G4013, G4014);
    or g_G4026 (G4026, G4015, G4016, G4017);
    or g_G4027 (G4027, G4018, G4019, G4020);
    or g_G4028 (G4028, G4021, G4022, G4023);
    or g_G4083 (G4083, G4070, G4071, G4072);
    or g_G4084 (G4084, G4073, G4074, G4075);
    or g_G4085 (G4085, G4076, G4077, G4078);
    or g_G4086 (G4086, G4079, G4080, G4081);
    nand g_G4368 (G4368, G4366, G4367);
    nand g_G4426 (G4426, G4424, G4425);
    not g_G4490 (G4490, G4484);
    nand g_G4493 (G4493, G4484, G4491);
    not g_G4578 (G4578, G4572);
    nand g_G4581 (G4581, G4572, G4579);
    nand g_G4832 (G4832, G4830, G4831);
    nand g_G4890 (G4890, G4888, G4889);
    nand g_G4948 (G4948, G4946, G4947);
    not g_G5032 (G5032, G5026);
    nand g_G5035 (G5035, G5026, G5033);
    and g_G642 (G642, G640, G1526);
    and g_G664 (G664, G662, G1606);
    and g_G667 (G667, G665, G1606);
    and g_G670 (G670, G668, G1606);
    and g_G676 (G676, G674, G2202);
    and g_G696 (G696, G694, G2279);
    and g_G699 (G699, G697, G2279);
    and g_G702 (G702, G700, G2279);
    and g_G811 (G811, G4113, G4096);
    and g_G812 (G812, G4096, G1936);
    and g_G818 (G818, G816, G817);
    and g_G853 (G853, G562, G853_tmp);
    and g_G853_tmp (G853_tmp, G3540, G3545, G3535, G3970);
    and g_G878 (G878, G3777, G3745, G3765);
    nand g_G4492 (G4492, G4487, G4490);
    nand g_G4580 (G4580, G4575, G4578);
    nand g_G5034 (G5034, G5029, G5032);
    and g_G1582 (G1582, G4083, G1540, G1564);
    and g_G1584 (G1584, G4025, G1528, G1564);
    and g_G1588 (G1588, G4084, G1540, G1564);
    and g_G1590 (G1590, G4026, G1528, G1564);
    and g_G1594 (G1594, G4085, G1540, G1564);
    and g_G1596 (G1596, G4027, G1528, G1564);
    and g_G1600 (G1600, G4086, G1540, G1564);
    and g_G1602 (G1602, G4028, G1528, G1564);
    and g_G2256 (G2256, G4083, G2215, G2238);
    and g_G2258 (G2258, G4025, G2203, G2238);
    and g_G2262 (G2262, G4084, G2215, G2238);
    and g_G2264 (G2264, G4026, G2203, G2238);
    and g_G2268 (G2268, G4085, G2215, G2238);
    and g_G2270 (G2270, G4027, G2203, G2238);
    and g_G2274 (G2274, G4086, G2215, G2238);
    and g_G2276 (G2276, G4028, G2203, G2238);
    and g_G708 (G708, G4086, G3672, G3696);
    and g_G709 (G709, G4028, G3660, G3696);
    and g_G723 (G723, G4086, G3570, G3594);
    and g_G724 (G724, G4028, G3558, G3594);
    and g_G728 (G728, G4085, G3570, G3594);
    and g_G729 (G729, G4027, G3558, G3594);
    and g_G733 (G733, G4084, G3570, G3594);
    and g_G734 (G734, G4026, G3558, G3594);
    and g_G738 (G738, G4083, G3570, G3594);
    and g_G739 (G739, G4025, G3558, G3594);
    and g_G768 (G768, G4085, G3672, G3696);
    and g_G769 (G769, G4027, G3660, G3696);
    and g_G773 (G773, G4084, G3672, G3696);
    and g_G774 (G774, G4026, G3660, G3696);
    and g_G778 (G778, G4083, G3672, G3696);
    and g_G779 (G779, G4025, G3660, G3696);
    or g_G813 (G813, G811, G812);
    not g_G824 (G824, G4086);
    not g_G826 (G826, G4085);
    not g_G828 (G828, G4084);
    not g_G830 (G830, G4083);
    and g_G854 (G854, G852, G853, G245);
    not g_G863 (G863, G4028);
    not g_G865 (G865, G4027);
    not g_G867 (G867, G4026);
    not g_G869 (G869, G4025);
    not g_G4374 (G4374, G4368);
    nand g_G4377 (G4377, G4368, G4375);
    not g_G4432 (G4432, G4426);
    nand g_G4435 (G4435, G4426, G4433);
    nand g_G4494 (G4494, G4492, G4493);
    nand g_G4582 (G4582, G4580, G4581);
    not g_G4838 (G4838, G4832);
    nand g_G4841 (G4841, G4832, G4839);
    not g_G4896 (G4896, G4890);
    nand g_G4899 (G4899, G4890, G4897);
    not g_G4954 (G4954, G4948);
    nand g_G4957 (G4957, G4948, G4955);
    nand g_G5036 (G5036, G5034, G5035);
    or g_G643 (G643, G1582, G1584, G1585, G1586);
    or g_G646 (G646, G1588, G1590, G1591, G1592);
    or g_G649 (G649, G1594, G1596, G1597, G1598);
    or g_G652 (G652, G1600, G1602, G1603, G1604);
    or g_G677 (G677, G2256, G2258, G2259, G2260);
    or g_G680 (G680, G2262, G2264, G2265, G2266);
    or g_G683 (G683, G2268, G2270, G2271, G2272);
    or g_G686 (G686, G2274, G2276, G2277, G2278);
    or g_G712 (G712, G708, G709, G710, G711);
    or g_G727 (G727, G723, G724, G725, G726);
    or g_G732 (G732, G728, G729, G730, G731);
    or g_G737 (G737, G733, G734, G735, G736);
    or g_G742 (G742, G738, G739, G740, G741);
    or g_G772 (G772, G768, G769, G770, G771);
    or g_G777 (G777, G773, G774, G775, G776);
    or g_G782 (G782, G778, G779, G780, G781);
    nand g_G4376 (G4376, G4371, G4374);
    nand g_G4434 (G4434, G4429, G4432);
    nand g_G4840 (G4840, G4835, G4838);
    nand g_G4898 (G4898, G4893, G4896);
    nand g_G4956 (G4956, G4951, G4954);
    and g_G645 (G645, G643, G1526);
    and g_G648 (G648, G646, G1526);
    and g_G651 (G651, G649, G1526);
    and g_G654 (G654, G652, G1526);
    and g_G679 (G679, G677, G2202);
    and g_G682 (G682, G680, G2202);
    and g_G685 (G685, G683, G2202);
    and g_G688 (G688, G686, G2202);
    nand g_G4378 (G4378, G4376, G4377);
    nand g_G4436 (G4436, G4434, G4435);
    not g_G4500 (G4500, G4494);
    nand g_G4503 (G4503, G4494, G4501);
    not g_G4588 (G4588, G4582);
    nand g_G4591 (G4591, G4582, G4589);
    nand g_G4842 (G4842, G4840, G4841);
    nand g_G4900 (G4900, G4898, G4899);
    nand g_G4958 (G4958, G4956, G4957);
    not g_G5042 (G5042, G5036);
    nand g_G5045 (G5045, G5036, G5043);
    nand g_G4502 (G4502, G4497, G4500);
    nand g_G4590 (G4590, G4585, G4588);
    nand g_G5044 (G5044, G5039, G5042);
    not g_G4384 (G4384, G4378);
    nand g_G4387 (G4387, G4378, G4385);
    not g_G4442 (G4442, G4436);
    nand g_G4445 (G4445, G4436, G4443);
    nand g_G4504 (G4504, G4502, G4503);
    nand g_G4592 (G4592, G4590, G4591);
    not g_G4848 (G4848, G4842);
    nand g_G4851 (G4851, G4842, G4849);
    not g_G4906 (G4906, G4900);
    nand g_G4909 (G4909, G4900, G4907);
    not g_G4964 (G4964, G4958);
    nand g_G4967 (G4967, G4958, G4965);
    nand g_G5046 (G5046, G5044, G5045);
    nand g_G4386 (G4386, G4381, G4384);
    nand g_G4444 (G4444, G4439, G4442);
    nand g_G4850 (G4850, G4845, G4848);
    nand g_G4908 (G4908, G4903, G4906);
    nand g_G4966 (G4966, G4961, G4964);
    nand g_G4388 (G4388, G4386, G4387);
    nand g_G4446 (G4446, G4444, G4445);
    not g_G4510 (G4510, G4504);
    nand g_G4513 (G4513, G4504, G4511);
    not g_G4598 (G4598, G4592);
    nand g_G4601 (G4601, G4592, G4599);
    nand g_G4852 (G4852, G4850, G4851);
    nand g_G4910 (G4910, G4908, G4909);
    nand g_G4968 (G4968, G4966, G4967);
    not g_G5052 (G5052, G5046);
    nand g_G5055 (G5055, G5046, G5053);
    nand g_G4512 (G4512, G4507, G4510);
    nand g_G4600 (G4600, G4595, G4598);
    nand g_G5054 (G5054, G5049, G5052);
    not g_G4394 (G4394, G4388);
    nand g_G4397 (G4397, G4388, G4395);
    not g_G4452 (G4452, G4446);
    nand g_G4455 (G4455, G4446, G4453);
    nand g_G4514 (G4514, G4512, G4513);
    nand g_G4602 (G4602, G4600, G4601);
    not g_G4858 (G4858, G4852);
    nand g_G4861 (G4861, G4852, G4859);
    not g_G4916 (G4916, G4910);
    nand g_G4919 (G4919, G4910, G4917);
    not g_G4974 (G4974, G4968);
    nand g_G4977 (G4977, G4968, G4975);
    nand g_G5056 (G5056, G5054, G5055);
    nand g_G4396 (G4396, G4391, G4394);
    nand g_G4454 (G4454, G4449, G4452);
    nand g_G4860 (G4860, G4855, G4858);
    nand g_G4918 (G4918, G4913, G4916);
    nand g_G4976 (G4976, G4971, G4974);
    nand g_G4398 (G4398, G4396, G4397);
    nand g_G4456 (G4456, G4454, G4455);
    not g_G4520 (G4520, G4514);
    nand g_G4523 (G4523, G4514, G4521);
    not g_G4608 (G4608, G4602);
    nand g_G4611 (G4611, G4602, G4609);
    nand g_G4862 (G4862, G4860, G4861);
    nand g_G4920 (G4920, G4918, G4919);
    nand g_G4978 (G4978, G4976, G4977);
    not g_G5062 (G5062, G5056);
    nand g_G5065 (G5065, G5056, G5063);
    nand g_G4522 (G4522, G4517, G4520);
    nand g_G4610 (G4610, G4605, G4608);
    nand g_G5064 (G5064, G5059, G5062);
    not g_G4404 (G4404, G4398);
    nand g_G1488 (G1488, G4398, G4405);
    not g_G4462 (G4462, G4456);
    nand g_G1493 (G1493, G4456, G4463);
    not g_G4868 (G4868, G4862);
    nand g_G2165 (G2165, G4862, G4869);
    not g_G4926 (G4926, G4920);
    nand g_G2170 (G2170, G4920, G4927);
    nand g_G4524 (G4524, G4522, G4523);
    nand g_G4612 (G4612, G4610, G4611);
    not g_G4984 (G4984, G4978);
    nand g_G4987 (G4987, G4978, G4985);
    nand g_G5066 (G5066, G5064, G5065);
    nand g_G1487 (G1487, G4401, G4404);
    nand g_G1492 (G1492, G4459, G4462);
    nand g_G2164 (G2164, G4865, G4868);
    nand g_G2169 (G2169, G4923, G4926);
    nand g_G4986 (G4986, G4981, G4984);
    nand g_G1489 (G1489, G1487, G1488);
    nand g_G1494 (G1494, G1492, G1493);
    nand g_G2166 (G2166, G2164, G2165);
    nand g_G2171 (G2171, G2169, G2170);
    not g_G4530 (G4530, G4524);
    nand g_G4533 (G4533, G4524, G4531);
    not g_G4618 (G4618, G4612);
    nand g_G4543 (G4543, G4612, G4619);
    nand g_G4988 (G4988, G4986, G4987);
    not g_G5072 (G5072, G5066);
    nand g_G4997 (G4997, G5066, G5073);
    nand g_G4532 (G4532, G4527, G4530);
    nand g_G4542 (G4542, G4615, G4618);
    nand g_G4996 (G4996, G5069, G5072);
    and g_G1513 (G1513, G1494, G1462, G1502);
    and g_G1514 (G1514, G1489, G1458, G1502);
    and g_G1515 (G1515, G1494, G1483, G1497);
    and g_G1516 (G1516, G1489, G1486, G1497);
    not g_G4994 (G4994, G4988);
    nand g_G2184 (G2184, G4988, G4995);
    and g_G2190 (G2190, G2171, G2139, G2179);
    and g_G2191 (G2191, G2166, G2135, G2179);
    and g_G2192 (G2192, G2171, G2160, G2174);
    and g_G2193 (G2193, G2166, G2163, G2174);
    nand g_G4534 (G4534, G4532, G4533);
    nand g_G4544 (G4544, G4542, G4543);
    nand g_G4998 (G4998, G4996, G4997);
    nand g_G2183 (G2183, G4991, G4994);
    or g_G4620 (G4620, G1513, G1514, G1515, G1516);
    or g_G5074 (G5074, G2190, G2191, G2192, G2193);
    not g_G4540 (G4540, G4534);
    nand g_G1507 (G1507, G4534, G4541);
    not g_G4550 (G4550, G4544);
    nand g_G1510 (G1510, G4544, G4551);
    nand g_G2185 (G2185, G2183, G2184);
    not g_G5004 (G5004, G4998);
    nand g_G2187 (G2187, G4998, G5005);
    nand g_G1506 (G1506, G4537, G4540);
    nand g_G1509 (G1509, G4547, G4550);
    not g_G4626 (G4626, G4620);
    nand g_G2186 (G2186, G5001, G5004);
    and g_G2195 (G2195, G2174, G2185);
    not g_G5080 (G5080, G5074);
    nand g_G1508 (G1508, G1506, G1507);
    nand g_G1511 (G1511, G1509, G1510);
    nand g_G2188 (G2188, G2186, G2187);
    not g_G1512 (G1512, G1511);
    and g_G1518 (G1518, G1497, G1508);
    not g_G2189 (G2189, G2188);
    and g_G1517 (G1517, G1512, G1502);
    and g_G2194 (G2194, G2189, G2179);
    or g_G4623 (G4623, G1517, G1518);
    or g_G5077 (G5077, G2194, G2195);
    nand g_G1519 (G1519, G4623, G4626);
    not g_G4627 (G4627, G4623);
    nand g_G2196 (G2196, G5077, G5080);
    not g_G5081 (G5081, G5077);
    nand g_G1520 (G1520, G4620, G4627);
    nand g_G2197 (G2197, G5074, G5081);
    nand g_G1521 (G1521, G1519, G1520);
    nand g_G2198 (G2198, G2196, G2197);
    and g_G840 (G840, G2198, G3795, G3823);
    and g_G879 (G879, G1521, G3737, G3765);
    not g_G1524 (G1524, G1521);
    not g_G2201 (G2201, G2198);
    or g_G843 (G843, G839, G840, G841, G842);
    or g_G882 (G882, G878, G879, G880, G881);
    and g_G3649 (G3649, G1524, G3628);
    and g_G3652 (G3652, G2201, G3628);
    or g_G3657 (G3657, G3648, G3649);
    or g_G3658 (G3658, G3651, G3652);
    and g_G3636 (G3636, G3657, G3622);
    and g_G3639 (G3639, G3658, G3622);
    and g_G3642 (G3642, G3657, G3622);
    and g_G3645 (G3645, G3658, G3622);
    or g_G3653 (G3653, G3636, G3637);
    or g_G3654 (G3654, G3639, G3640);
    or g_G3655 (G3655, G3642, G3643);
    or g_G3656 (G3656, G3645, G3646);
    and g_G763 (G763, G3656, G2430, G2454);
    and g_G764 (G764, G3655, G2418, G2454);
    and g_G803 (G803, G3656, G2488, G2512);
    and g_G804 (G804, G3655, G2476, G2512);
    and g_G1657 (G1657, G3654, G1621, G1645);
    and g_G1659 (G1659, G3653, G1609, G1645);
    and g_G2328 (G2328, G3654, G2293, G2316);
    and g_G2330 (G2330, G3653, G2281, G2316);
    or g_G1662 (G1662, G1657, G1659, G1660, G1661);
    or g_G2333 (G2333, G2328, G2330, G2331, G2332);
    or g_G767 (G767, G763, G764, G765, G766);
    or g_G807 (G807, G803, G804, G805, G806);
    and g_G657 (G657, G1662, G1606);
    and g_G689 (G689, G2333, G2279);
    not g_G658 (G658, G657);
    not g_G690 (G690, G689);

endmodule
