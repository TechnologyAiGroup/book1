module s444(clk,G0,G1,G2,G118,G167,G107,G119,G168,G108);
	input clk,G0,G1,G2;
    output G118,G167,G107,G119,G168,G108;

	sky130_fd_sc_hd__dfxtp_1 g_G11 ( .D(G37), .CLK(clk), .Q(G11) );
	sky130_fd_sc_hd__dfxtp_1 g_G12 ( .D(G41), .CLK(clk), .Q(G12) );
	sky130_fd_sc_hd__dfxtp_1 g_G13 ( .D(G45), .CLK(clk), .Q(G13) );
	sky130_fd_sc_hd__dfxtp_1 g_G14 ( .D(G49), .CLK(clk), .Q(G14) );
	sky130_fd_sc_hd__dfxtp_1 g_G15 ( .D(G58), .CLK(clk), .Q(G15) );
    sky130_fd_sc_hd__dfxtp_1 g_G16 ( .D(G62), .CLK(clk), .Q(G16) );
	sky130_fd_sc_hd__dfxtp_1 g_G17 ( .D(G66), .CLK(clk), .Q(G17) );
	sky130_fd_sc_hd__dfxtp_1 g_G18 ( .D(G70), .CLK(clk), .Q(G18) );
	sky130_fd_sc_hd__dfxtp_1 g_G19 ( .D(G80), .CLK(clk), .Q(G19) );
	sky130_fd_sc_hd__dfxtp_1 g_G20 ( .D(G84), .CLK(clk), .Q(G20) );
	sky130_fd_sc_hd__dfxtp_1 g_G21 ( .D(G88), .CLK(clk), .Q(G21) );
	sky130_fd_sc_hd__dfxtp_1 g_G22 ( .D(G92), .CLK(clk), .Q(G22) );
	sky130_fd_sc_hd__dfxtp_1 g_G23 ( .D(G101), .CLK(clk), .Q(G23) );
	sky130_fd_sc_hd__dfxtp_1 g_G24 ( .D(G162BF), .CLK(clk), .Q(G24) );
	sky130_fd_sc_hd__dfxtp_1 g_G25 ( .D(G109), .CLK(clk), .Q(G25) );
	sky130_fd_sc_hd__dfxtp_1 g_G26 ( .D(G110), .CLK(clk), .Q(G26) );
	sky130_fd_sc_hd__dfxtp_1 g_G27 ( .D(G111), .CLK(clk), .Q(G27) );
	sky130_fd_sc_hd__dfxtp_1 g_G28 ( .D(G112), .CLK(clk), .Q(G28) );
	sky130_fd_sc_hd__dfxtp_1 g_G29 ( .D(G113), .CLK(clk), .Q(G29) );
	sky130_fd_sc_hd__dfxtp_1 g_G30 ( .D(G114), .CLK(clk), .Q(G30) );
	sky130_fd_sc_hd__dfxtp_1 g_G31 ( .D(G155), .CLK(clk), .Q(G31) );
	sky130_fd_sc_hd__inv_1 g_I372 ( .A(G0), .Y(I372) );
	sky130_fd_sc_hd__inv_1 g_I382 ( .A(G1), .Y(I382) );
	sky130_fd_sc_hd__inv_1 g_I318 ( .A(G2), .Y(I318) );
	sky130_fd_sc_hd__inv_1 g_G34 ( .A(G11), .Y(G34) );
	sky130_fd_sc_hd__inv_1 g_I180 ( .A(G11), .Y(I180) );
	sky130_fd_sc_hd__inv_1 g_G35 ( .A(G12), .Y(G35) );
	sky130_fd_sc_hd__inv_1 g_G77 ( .A(G20), .Y(G77) );
	sky130_fd_sc_hd__inv_1 g_G135 ( .A(G20), .Y(G135) );
	sky130_fd_sc_hd__inv_1 g_G36 ( .A(G13), .Y(G36) );
	sky130_fd_sc_hd__inv_1 g_G78 ( .A(G21), .Y(G78) );
	sky130_fd_sc_hd__inv_1 g_G144 ( .A(G21), .Y(G144) );
	sky130_fd_sc_hd__inv_1 g_G32 ( .A(G14), .Y(G32) );
	sky130_fd_sc_hd__inv_1 g_G74 ( .A(G22), .Y(G74) );
	sky130_fd_sc_hd__inv_1 g_G142 ( .A(G22), .Y(G142) );
	sky130_fd_sc_hd__inv_1 g_I392 ( .A(G30), .Y(I392) );
	sky130_fd_sc_hd__inv_1 g_G55 ( .A(G15), .Y(G55) );
	sky130_fd_sc_hd__inv_1 g_G102 ( .A(G23), .Y(G102) );
	sky130_fd_sc_hd__inv_1 g_G136 ( .A(G23), .Y(G136) );
	sky130_fd_sc_hd__inv_1 g_G156 ( .A(G31), .Y(G156) );
	sky130_fd_sc_hd__inv_1 g_G56 ( .A(G16), .Y(G56) );
	sky130_fd_sc_hd__inv_1 g_G143 ( .A(G24), .Y(G143) );
	sky130_fd_sc_hd__inv_1 g_G161 ( .A(G17), .Y(G161) );
	sky130_fd_sc_hd__inv_1 g_I321 ( .A(G25), .Y(I321) );
	sky130_fd_sc_hd__inv_1 g_G53 ( .A(G18), .Y(G53) );
	sky130_fd_sc_hd__inv_1 g_I324 ( .A(G26), .Y(I324) );
	sky130_fd_sc_hd__inv_1 g_G76 ( .A(G19), .Y(G76) );
	sky130_fd_sc_hd__inv_1 g_G150 ( .A(G19), .Y(G150) );
	sky130_fd_sc_hd__inv_1 g_I336 ( .A(G27), .Y(I336) );
	sky130_fd_sc_hd__inv_1 g_G119 ( .A(G28), .Y(G119) );
	sky130_fd_sc_hd__inv_1 g_G167 ( .A(G29), .Y(G167) );
	sky130_fd_sc_hd__inv_1 g_G152 ( .A(I372), .Y(G152) );
	sky130_fd_sc_hd__inv_1 g_G160 ( .A(I382), .Y(G160) );
	sky130_fd_sc_hd__inv_1 g_G106 ( .A(I318), .Y(G106) );
	sky130_fd_sc_hd__inv_1 g_G43 ( .A(G34), .Y(G43) );
	sky130_fd_sc_hd__inv_1 g_I182 ( .A(I180), .Y(I182) );
	sky130_fd_sc_hd__inv_1 g_G168 ( .A(I392), .Y(G168) );
	sky130_fd_sc_hd__inv_1 g_G107 ( .A(I321), .Y(G107) );
	sky130_fd_sc_hd__inv_1 g_G108 ( .A(I324), .Y(G108) );
	sky130_fd_sc_hd__inv_1 g_G118 ( .A(I336), .Y(G118) );
	sky130_fd_sc_hd__inv_1 g_G99 ( .A(G152), .Y(G99) );
	sky130_fd_sc_hd__inv_1 g_G139 ( .A(G152), .Y(G139) );
	sky130_fd_sc_hd__inv_1 g_G153 ( .A(G152), .Y(G153) );
	sky130_fd_sc_hd__inv_1 g_G157 ( .A(G160), .Y(G157) );
	sky130_fd_sc_hd__inv_1 g_G103 ( .A(G106), .Y(G103) );
	sky130_fd_sc_hd__inv_1 g_G38 ( .A(G40), .Y(G38) );
	sky130_fd_sc_hd__inv_1 g_G60 ( .A(G57), .Y(G60) );
	sky130_fd_sc_hd__inv_1 g_G79 ( .A(G97), .Y(G79) );
	sky130_fd_sc_hd__inv_1 g_G42 ( .A(G44), .Y(G42) );
	sky130_fd_sc_hd__inv_1 g_G46 ( .A(G48), .Y(G46) );
	sky130_fd_sc_hd__inv_1 g_I105 ( .A(G162), .Y(I105) );
	sky130_fd_sc_hd__inv_1 g_G166 ( .A(G162), .Y(G166) );
	sky130_fd_sc_hd__inv_1 g_G50 ( .A(G52), .Y(G50) );
	sky130_fd_sc_hd__inv_1 g_G82 ( .A(G79), .Y(G82) );
	sky130_fd_sc_hd__inv_1 g_G162BF ( .A(I105), .Y(G162BF) );
	sky130_fd_sc_hd__inv_1 g_G59 ( .A(G61), .Y(G59) );
	sky130_fd_sc_hd__inv_1 g_G63 ( .A(G65), .Y(G63) );
	sky130_fd_sc_hd__inv_1 g_G67 ( .A(G69), .Y(G67) );
	sky130_fd_sc_hd__inv_1 g_G71 ( .A(G73), .Y(G71) );
	sky130_fd_sc_hd__inv_1 g_G81 ( .A(G83), .Y(G81) );
	sky130_fd_sc_hd__inv_1 g_G85 ( .A(G87), .Y(G85) );
	sky130_fd_sc_hd__inv_1 g_G89 ( .A(G91), .Y(G89) );
	sky130_fd_sc_hd__inv_1 g_G94 ( .A(G96), .Y(G94) );
	sky130_fd_sc_hd__and2_1 g_G122 ( .A(G24), .B(G121), .X(G122) );
	sky130_fd_sc_hd__and3_1 g_G124 ( .A(G139), .B(G22), .C(G150), .X(G124) );
	sky130_fd_sc_hd__and3_1 g_G125 ( .A(G139), .B(G20), .C(G19), .X(G125) );
	sky130_fd_sc_hd__and2_1 g_G126 ( .A(G139), .B(G21), .X(G126) );
	sky130_fd_sc_hd__and2_1 g_G127 ( .A(G139), .B(G24), .X(G127) );
	sky130_fd_sc_hd__and2_1 g_G154 ( .A(G158), .B(G159), .X(G154) );
	sky130_fd_sc_hd__and2_1 g_G100 ( .A(G104), .B(G105), .X(G100) );
	sky130_fd_sc_hd__and2_1 g_G155 ( .A(G154), .B(G153), .X(G155) );
	sky130_fd_sc_hd__and2_1 g_G101 ( .A(G100), .B(G99), .X(G101) );
	sky130_fd_sc_hd__and3_1 g_G115 ( .A(G161), .B(G117), .C(G162), .X(G115) );
	sky130_fd_sc_hd__and3_1 g_G163 ( .A(G161), .B(G165), .C(G162), .X(G163) );
	sky130_fd_sc_hd__and2_1 g_G116 ( .A(G117), .B(G166), .X(G116) );
	sky130_fd_sc_hd__and2_1 g_G164 ( .A(G165), .B(G166), .X(G164) );
	sky130_fd_sc_hd__or3_1 g_G141 ( .A(G24), .B(G22), .C(G21), .X(G141) );
	sky130_fd_sc_hd__or3_1 g_G137 ( .A(G136), .B(G20), .C(G19), .X(G137) );
	sky130_fd_sc_hd__or2_1 g_G138 ( .A(G136), .B(G142), .X(G138) );
	sky130_fd_sc_hd__or4_1 g_G140 ( .A(G24), .B(G21), .C(G20), .D(G150), .X(G140) );
	sky130_fd_sc_hd__or4_1 g_G133 ( .A(G152), .B(G136), .C(G22), .D(G144), .X(G133) );
	sky130_fd_sc_hd__or3_1 g_G134 ( .A(G152), .B(G142), .C(G21), .X(G134) );
	sky130_fd_sc_hd__or4_1 g_G145 ( .A(G152), .B(G142), .C(G20), .D(G19), .X(G145) );
	sky130_fd_sc_hd__or2_1 g_G146 ( .A(G152), .B(G143), .X(G146) );
	sky130_fd_sc_hd__or2_1 g_G147 ( .A(G152), .B(G144), .X(G147) );
	sky130_fd_sc_hd__or2_1 g_G158 ( .A(G31), .B(G160), .X(G158) );
	sky130_fd_sc_hd__or2_1 g_G104 ( .A(G23), .B(G106), .X(G104) );
	sky130_fd_sc_hd__or4_1 g_G131 ( .A(G144), .B(G22), .C(G23), .D(G129), .X(G131) );
	sky130_fd_sc_hd__or2_1 g_G159 ( .A(G156), .B(G157), .X(G159) );
	sky130_fd_sc_hd__or2_1 g_G105 ( .A(G102), .B(G103), .X(G105) );
	sky130_fd_sc_hd__nand2_1 g_I181 ( .A(G11), .B(I180), .Y(I181) );
	sky130_fd_sc_hd__nand2_1 g_G129 ( .A(G19), .B(G135), .Y(G129) );
	sky130_fd_sc_hd__nand4_1 g_G121 ( .A(G19), .B(G135), .C(G142), .D(G136), .Y(G121) );
	sky130_fd_sc_hd__nand2_1 g_I190 ( .A(G12), .B(G43), .Y(I190) );
	sky130_fd_sc_hd__nand2_1 g_G40 ( .A(I181), .B(I182), .Y(G40) );
	sky130_fd_sc_hd__nand2_1 g_I200 ( .A(G13), .B(G47), .Y(I200) );
	sky130_fd_sc_hd__nand2_1 g_I210 ( .A(G14), .B(G51), .Y(I210) );
	sky130_fd_sc_hd__nand2_1 g_G120 ( .A(G150), .B(G128), .Y(G120) );
	sky130_fd_sc_hd__nand2_1 g_G132 ( .A(G133), .B(G134), .Y(G132) );
	sky130_fd_sc_hd__nand3_1 g_G111 ( .A(G140), .B(G141), .C(G139), .Y(G111) );
	sky130_fd_sc_hd__nand4_1 g_G123 ( .A(G137), .B(G138), .C(G21), .D(G139), .Y(G123) );
	sky130_fd_sc_hd__nand4_1 g_G151 ( .A(G20), .B(G144), .C(G143), .D(G139), .Y(G151) );
	sky130_fd_sc_hd__nand3_1 g_G117 ( .A(G145), .B(G146), .C(G147), .Y(G117) );
	sky130_fd_sc_hd__nand2_1 g_I191 ( .A(G12), .B(I190), .Y(I191) );
	sky130_fd_sc_hd__nand2_1 g_I192 ( .A(G43), .B(I190), .Y(I192) );
	sky130_fd_sc_hd__nand2_1 g_I201 ( .A(G13), .B(I200), .Y(I201) );
	sky130_fd_sc_hd__nand2_1 g_I202 ( .A(G47), .B(I200), .Y(I202) );
	sky130_fd_sc_hd__nand2_1 g_G149 ( .A(G131), .B(G130), .Y(G149) );
	sky130_fd_sc_hd__nand2_1 g_I211 ( .A(G14), .B(I210), .Y(I211) );
	sky130_fd_sc_hd__nand2_1 g_I212 ( .A(G51), .B(I210), .Y(I212) );
	sky130_fd_sc_hd__nand3_1 g_G148 ( .A(G150), .B(G135), .C(G132), .Y(G148) );
	sky130_fd_sc_hd__nand2_1 g_G44 ( .A(I191), .B(I192), .Y(G44) );
	sky130_fd_sc_hd__nand2_1 g_G48 ( .A(I201), .B(I202), .Y(G48) );
	sky130_fd_sc_hd__nand2_1 g_G162 ( .A(G120), .B(G149), .Y(G162) );
	sky130_fd_sc_hd__nand2_1 g_G52 ( .A(I211), .B(I212), .Y(G52) );
	sky130_fd_sc_hd__nand2_1 g_I225 ( .A(G15), .B(G60), .Y(I225) );
	sky130_fd_sc_hd__nand2_1 g_I235 ( .A(G16), .B(G64), .Y(I235) );
	sky130_fd_sc_hd__nand2_1 g_I245 ( .A(G17), .B(G68), .Y(I245) );
	sky130_fd_sc_hd__nand2_1 g_I255 ( .A(G18), .B(G72), .Y(I255) );
	sky130_fd_sc_hd__nand2_1 g_G165 ( .A(G148), .B(G149), .Y(G165) );
	sky130_fd_sc_hd__nand2_1 g_I226 ( .A(G15), .B(I225), .Y(I226) );
	sky130_fd_sc_hd__nand2_1 g_I227 ( .A(G60), .B(I225), .Y(I227) );
	sky130_fd_sc_hd__nand2_1 g_I236 ( .A(G16), .B(I235), .Y(I236) );
	sky130_fd_sc_hd__nand2_1 g_I237 ( .A(G64), .B(I235), .Y(I237) );
	sky130_fd_sc_hd__nand2_1 g_I246 ( .A(G17), .B(I245), .Y(I246) );
	sky130_fd_sc_hd__nand2_1 g_I247 ( .A(G68), .B(I245), .Y(I247) );
	sky130_fd_sc_hd__nand2_1 g_I256 ( .A(G18), .B(I255), .Y(I256) );
	sky130_fd_sc_hd__nand2_1 g_I257 ( .A(G72), .B(I255), .Y(I257) );
	sky130_fd_sc_hd__nand2_1 g_G61 ( .A(I226), .B(I227), .Y(G61) );
	sky130_fd_sc_hd__nand2_1 g_G65 ( .A(I236), .B(I237), .Y(G65) );
	sky130_fd_sc_hd__nand2_1 g_G69 ( .A(I246), .B(I247), .Y(G69) );
	sky130_fd_sc_hd__nand2_1 g_G73 ( .A(I256), .B(I257), .Y(G73) );
	sky130_fd_sc_hd__nand2_1 g_I271 ( .A(G19), .B(G82), .Y(I271) );
	sky130_fd_sc_hd__nand2_1 g_I281 ( .A(G20), .B(G86), .Y(I281) );
	sky130_fd_sc_hd__nand2_1 g_I291 ( .A(G21), .B(G90), .Y(I291) );
	sky130_fd_sc_hd__nand2_1 g_I302 ( .A(G22), .B(G95), .Y(I302) );
	sky130_fd_sc_hd__nand2_1 g_I272 ( .A(G19), .B(I271), .Y(I272) );
	sky130_fd_sc_hd__nand2_1 g_I273 ( .A(G82), .B(I271), .Y(I273) );
	sky130_fd_sc_hd__nand2_1 g_I282 ( .A(G20), .B(I281), .Y(I282) );
	sky130_fd_sc_hd__nand2_1 g_I283 ( .A(G86), .B(I281), .Y(I283) );
	sky130_fd_sc_hd__nand2_1 g_I292 ( .A(G21), .B(I291), .Y(I292) );
	sky130_fd_sc_hd__nand2_1 g_I293 ( .A(G90), .B(I291), .Y(I293) );
	sky130_fd_sc_hd__nand2_1 g_I303 ( .A(G22), .B(I302), .Y(I303) );
	sky130_fd_sc_hd__nand2_1 g_I304 ( .A(G95), .B(I302), .Y(I304) );
	sky130_fd_sc_hd__nand2_1 g_G83 ( .A(I272), .B(I273), .Y(G83) );
	sky130_fd_sc_hd__nand2_1 g_G87 ( .A(I282), .B(I283), .Y(G87) );
	sky130_fd_sc_hd__nand2_1 g_G91 ( .A(I292), .B(I293), .Y(G91) );
	sky130_fd_sc_hd__nand2_1 g_G96 ( .A(I303), .B(I304), .Y(G96) );
	sky130_fd_sc_hd__nor3_1 g_G33 ( .A(G11), .B(G12), .C(G13), .Y(G33) );
	sky130_fd_sc_hd__nor3_1 g_G54 ( .A(G15), .B(G16), .C(G17), .Y(G54) );
	sky130_fd_sc_hd__nor3_1 g_G75 ( .A(G19), .B(G20), .C(G21), .Y(G75) );
	sky130_fd_sc_hd__nor2_1 g_G47 ( .A(G34), .B(G35), .Y(G47) );
	sky130_fd_sc_hd__nor3_1 g_G51 ( .A(G34), .B(G35), .C(G36), .Y(G51) );
	sky130_fd_sc_hd__nor2_1 g_G98 ( .A(G32), .B(G33), .Y(G98) );
	sky130_fd_sc_hd__nor4_1 g_G128 ( .A(G20), .B(G144), .C(G136), .D(G152), .Y(G128) );
	sky130_fd_sc_hd__nor2_1 g_G130 ( .A(G143), .B(G152), .Y(G130) );
	sky130_fd_sc_hd__nor2_1 g_G57 ( .A(G31), .B(G98), .Y(G57) );
	sky130_fd_sc_hd__nor2_1 g_G64 ( .A(G55), .B(G57), .Y(G64) );
	sky130_fd_sc_hd__nor3_1 g_G68 ( .A(G55), .B(G56), .C(G57), .Y(G68) );
	sky130_fd_sc_hd__nor4_1 g_G72 ( .A(G55), .B(G56), .C(G161), .D(G57), .Y(G72) );
	sky130_fd_sc_hd__nor3_1 g_G97 ( .A(G53), .B(G57), .C(G54), .Y(G97) );
	sky130_fd_sc_hd__nor2_1 g_G109 ( .A(G122), .B(G123), .Y(G109) );
	sky130_fd_sc_hd__nor4_1 g_G110 ( .A(G124), .B(G125), .C(G126), .D(G127), .Y(G110) );
	sky130_fd_sc_hd__nor2_1 g_G114 ( .A(G150), .B(G151), .Y(G114) );
	sky130_fd_sc_hd__nor3_1 g_G37 ( .A(G98), .B(G38), .C(G152), .Y(G37) );
	sky130_fd_sc_hd__nor2_1 g_G86 ( .A(G76), .B(G79), .Y(G86) );
	sky130_fd_sc_hd__nor3_1 g_G90 ( .A(G76), .B(G77), .C(G79), .Y(G90) );
	sky130_fd_sc_hd__nor3_1 g_G93 ( .A(G74), .B(G79), .C(G75), .Y(G93) );
	sky130_fd_sc_hd__nor4_1 g_G95 ( .A(G76), .B(G77), .C(G78), .D(G79), .Y(G95) );
	sky130_fd_sc_hd__nor3_1 g_G41 ( .A(G98), .B(G42), .C(G152), .Y(G41) );
	sky130_fd_sc_hd__nor3_1 g_G45 ( .A(G98), .B(G46), .C(G152), .Y(G45) );
	sky130_fd_sc_hd__nor3_1 g_G49 ( .A(G98), .B(G50), .C(G152), .Y(G49) );
	sky130_fd_sc_hd__nor2_1 g_G112 ( .A(G115), .B(G116), .Y(G112) );
	sky130_fd_sc_hd__nor2_1 g_G113 ( .A(G163), .B(G164), .Y(G113) );
	sky130_fd_sc_hd__nor3_1 g_G58 ( .A(G97), .B(G59), .C(G152), .Y(G58) );
	sky130_fd_sc_hd__nor3_1 g_G62 ( .A(G97), .B(G63), .C(G152), .Y(G62) );
	sky130_fd_sc_hd__nor3_1 g_G66 ( .A(G97), .B(G67), .C(G152), .Y(G66) );
	sky130_fd_sc_hd__nor3_1 g_G70 ( .A(G97), .B(G71), .C(G152), .Y(G70) );
	sky130_fd_sc_hd__nor3_1 g_G80 ( .A(G93), .B(G81), .C(G152), .Y(G80) );
	sky130_fd_sc_hd__nor3_1 g_G84 ( .A(G93), .B(G85), .C(G152), .Y(G84) );
	sky130_fd_sc_hd__nor3_1 g_G88 ( .A(G93), .B(G89), .C(G152), .Y(G88) );
	sky130_fd_sc_hd__nor3_1 g_G92 ( .A(G93), .B(G94), .C(G152), .Y(G92) );
	
endmodule
		